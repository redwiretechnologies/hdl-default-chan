// SPDX-License-Identifier: Apache-2.0

/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : pfb_128Mmax_16iw_16ow_32tps_dp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data
//
//
/*****************************************************************************/


module pfb_128Mmax_16iw_16ow_32tps_dp_rom
(
  input clk,
  input wea,
  input [24:0] dia,
  input [11:0] addra,
  input [11:0] addrb,
  output [24:0] dob
);

(* rom_style = "block" *) reg [24:0] rom [4095:0];
reg [11:0] addrb_d;
reg [24:0] dob_d;
reg [24:0] rom_pipea;
reg [11:0] addra_d;
reg [24:0] dia_d;
reg wea_d;

assign dob = dob_d;

initial
begin
    rom[0] = 25'b1111111111111111000001011;
    rom[1] = 25'b1111111111111111000001011;
    rom[2] = 25'b1111111111111111000001010;
    rom[3] = 25'b1111111111111111000001010;
    rom[4] = 25'b1111111111111111000001000;
    rom[5] = 25'b1111111111111111000000111;
    rom[6] = 25'b1111111111111111000000100;
    rom[7] = 25'b1111111111111111000000010;
    rom[8] = 25'b1111111111111111000000000;
    rom[9] = 25'b1111111111111110111111101;
    rom[10] = 25'b1111111111111110111111001;
    rom[11] = 25'b1111111111111110111110110;
    rom[12] = 25'b1111111111111110111110010;
    rom[13] = 25'b1111111111111110111101101;
    rom[14] = 25'b1111111111111110111101001;
    rom[15] = 25'b1111111111111110111100100;
    rom[16] = 25'b1111111111111110111011110;
    rom[17] = 25'b1111111111111110111011001;
    rom[18] = 25'b1111111111111110111010011;
    rom[19] = 25'b1111111111111110111001100;
    rom[20] = 25'b1111111111111110111000111;
    rom[21] = 25'b1111111111111110110111111;
    rom[22] = 25'b1111111111111110110111000;
    rom[23] = 25'b1111111111111110110110001;
    rom[24] = 25'b1111111111111110110101001;
    rom[25] = 25'b1111111111111110110100001;
    rom[26] = 25'b1111111111111110110011001;
    rom[27] = 25'b1111111111111110110010000;
    rom[28] = 25'b1111111111111110110001000;
    rom[29] = 25'b1111111111111110101111111;
    rom[30] = 25'b1111111111111110101110101;
    rom[31] = 25'b1111111111111110101101100;
    rom[32] = 25'b1111111111111110101100011;
    rom[33] = 25'b1111111111111110101011000;
    rom[34] = 25'b1111111111111110101001110;
    rom[35] = 25'b1111111111111110101000100;
    rom[36] = 25'b1111111111111110100111010;
    rom[37] = 25'b1111111111111110100101110;
    rom[38] = 25'b1111111111111110100100100;
    rom[39] = 25'b1111111111111110100011001;
    rom[40] = 25'b1111111111111110100001110;
    rom[41] = 25'b1111111111111110100000010;
    rom[42] = 25'b1111111111111110011110111;
    rom[43] = 25'b1111111111111110011101011;
    rom[44] = 25'b1111111111111110011100000;
    rom[45] = 25'b1111111111111110011010100;
    rom[46] = 25'b1111111111111110011001000;
    rom[47] = 25'b1111111111111110010111100;
    rom[48] = 25'b1111111111111110010110000;
    rom[49] = 25'b1111111111111110010100100;
    rom[50] = 25'b1111111111111110010011000;
    rom[51] = 25'b1111111111111110010001101;
    rom[52] = 25'b1111111111111110010000001;
    rom[53] = 25'b1111111111111110001110100;
    rom[54] = 25'b1111111111111110001101000;
    rom[55] = 25'b1111111111111110001011100;
    rom[56] = 25'b1111111111111110001010000;
    rom[57] = 25'b1111111111111110001000100;
    rom[58] = 25'b1111111111111110000111000;
    rom[59] = 25'b1111111111111110000101100;
    rom[60] = 25'b1111111111111110000100000;
    rom[61] = 25'b1111111111111110000010100;
    rom[62] = 25'b1111111111111110000001001;
    rom[63] = 25'b1111111111111101111111101;
    rom[64] = 25'b1111111111111101111110010;
    rom[65] = 25'b1111111111111101111100111;
    rom[66] = 25'b1111111111111101111011101;
    rom[67] = 25'b1111111111111101111010001;
    rom[68] = 25'b1111111111111101111000111;
    rom[69] = 25'b1111111111111101110111100;
    rom[70] = 25'b1111111111111101110110010;
    rom[71] = 25'b1111111111111101110101000;
    rom[72] = 25'b1111111111111101110011110;
    rom[73] = 25'b1111111111111101110010100;
    rom[74] = 25'b1111111111111101110001011;
    rom[75] = 25'b1111111111111101110000010;
    rom[76] = 25'b1111111111111101101111001;
    rom[77] = 25'b1111111111111101101110001;
    rom[78] = 25'b1111111111111101101101001;
    rom[79] = 25'b1111111111111101101100010;
    rom[80] = 25'b1111111111111101101011010;
    rom[81] = 25'b1111111111111101101010011;
    rom[82] = 25'b1111111111111101101001100;
    rom[83] = 25'b1111111111111101101000110;
    rom[84] = 25'b1111111111111101101000000;
    rom[85] = 25'b1111111111111101100111011;
    rom[86] = 25'b1111111111111101100110110;
    rom[87] = 25'b1111111111111101100110000;
    rom[88] = 25'b1111111111111101100101101;
    rom[89] = 25'b1111111111111101100101001;
    rom[90] = 25'b1111111111111101100100101;
    rom[91] = 25'b1111111111111101100100011;
    rom[92] = 25'b1111111111111101100100001;
    rom[93] = 25'b1111111111111101100011110;
    rom[94] = 25'b1111111111111101100011101;
    rom[95] = 25'b1111111111111101100011100;
    rom[96] = 25'b1111111111111101100011100;
    rom[97] = 25'b1111111111111101100011100;
    rom[98] = 25'b1111111111111101100011110;
    rom[99] = 25'b1111111111111101100011111;
    rom[100] = 25'b1111111111111101100100001;
    rom[101] = 25'b1111111111111101100100100;
    rom[102] = 25'b1111111111111101100100111;
    rom[103] = 25'b1111111111111101100101010;
    rom[104] = 25'b1111111111111101100101111;
    rom[105] = 25'b1111111111111101100110100;
    rom[106] = 25'b1111111111111101100111010;
    rom[107] = 25'b1111111111111101101000001;
    rom[108] = 25'b1111111111111101101000111;
    rom[109] = 25'b1111111111111101101001111;
    rom[110] = 25'b1111111111111101101011000;
    rom[111] = 25'b1111111111111101101100001;
    rom[112] = 25'b1111111111111101101101010;
    rom[113] = 25'b1111111111111101101110101;
    rom[114] = 25'b1111111111111101110000000;
    rom[115] = 25'b1111111111111101110001100;
    rom[116] = 25'b1111111111111101110011001;
    rom[117] = 25'b1111111111111101110100110;
    rom[118] = 25'b1111111111111101110110100;
    rom[119] = 25'b1111111111111101111000011;
    rom[120] = 25'b1111111111111101111010011;
    rom[121] = 25'b1111111111111101111100011;
    rom[122] = 25'b1111111111111101111110100;
    rom[123] = 25'b1111111111111110000000110;
    rom[124] = 25'b1111111111111110000011000;
    rom[125] = 25'b1111111111111110000101100;
    rom[126] = 25'b1111111111111110001000000;
    rom[127] = 25'b1111111111111110001010101;
    rom[128] = 25'b1111111111111110001101011;
    rom[129] = 25'b1111111111111110010000001;
    rom[130] = 25'b1111111111111110010011000;
    rom[131] = 25'b1111111111111110010110000;
    rom[132] = 25'b1111111111111110011001010;
    rom[133] = 25'b1111111111111110011100011;
    rom[134] = 25'b1111111111111110011111101;
    rom[135] = 25'b1111111111111110100011001;
    rom[136] = 25'b1111111111111110100110100;
    rom[137] = 25'b1111111111111110101010001;
    rom[138] = 25'b1111111111111110101101111;
    rom[139] = 25'b1111111111111110110001101;
    rom[140] = 25'b1111111111111110110101100;
    rom[141] = 25'b1111111111111110111001100;
    rom[142] = 25'b1111111111111110111101101;
    rom[143] = 25'b1111111111111111000001111;
    rom[144] = 25'b1111111111111111000110001;
    rom[145] = 25'b1111111111111111001010011;
    rom[146] = 25'b1111111111111111001110111;
    rom[147] = 25'b1111111111111111010011100;
    rom[148] = 25'b1111111111111111011000001;
    rom[149] = 25'b1111111111111111011100111;
    rom[150] = 25'b1111111111111111100001110;
    rom[151] = 25'b1111111111111111100110101;
    rom[152] = 25'b1111111111111111101011110;
    rom[153] = 25'b1111111111111111110000111;
    rom[154] = 25'b1111111111111111110110000;
    rom[155] = 25'b1111111111111111111011011;
    rom[156] = 25'b0000000000000000000000101;
    rom[157] = 25'b0000000000000000000110001;
    rom[158] = 25'b0000000000000000001011101;
    rom[159] = 25'b0000000000000000010001011;
    rom[160] = 25'b0000000000000000010111000;
    rom[161] = 25'b0000000000000000011100111;
    rom[162] = 25'b0000000000000000100010110;
    rom[163] = 25'b0000000000000000101000101;
    rom[164] = 25'b0000000000000000101110110;
    rom[165] = 25'b0000000000000000110100111;
    rom[166] = 25'b0000000000000000111011000;
    rom[167] = 25'b0000000000000001000001010;
    rom[168] = 25'b0000000000000001000111101;
    rom[169] = 25'b0000000000000001001110000;
    rom[170] = 25'b0000000000000001010100100;
    rom[171] = 25'b0000000000000001011011000;
    rom[172] = 25'b0000000000000001100001101;
    rom[173] = 25'b0000000000000001101000010;
    rom[174] = 25'b0000000000000001101111000;
    rom[175] = 25'b0000000000000001110101110;
    rom[176] = 25'b0000000000000001111100101;
    rom[177] = 25'b0000000000000010000011100;
    rom[178] = 25'b0000000000000010001010100;
    rom[179] = 25'b0000000000000010010001011;
    rom[180] = 25'b0000000000000010011000100;
    rom[181] = 25'b0000000000000010011111100;
    rom[182] = 25'b0000000000000010100110101;
    rom[183] = 25'b0000000000000010101101110;
    rom[184] = 25'b0000000000000010110101000;
    rom[185] = 25'b0000000000000010111100001;
    rom[186] = 25'b0000000000000011000011011;
    rom[187] = 25'b0000000000000011001010101;
    rom[188] = 25'b0000000000000011010010000;
    rom[189] = 25'b0000000000000011011001011;
    rom[190] = 25'b0000000000000011100000101;
    rom[191] = 25'b0000000000000011101000000;
    rom[192] = 25'b0000000000000011101111011;
    rom[193] = 25'b0000000000000011110110110;
    rom[194] = 25'b0000000000000011111110010;
    rom[195] = 25'b0000000000000100000101101;
    rom[196] = 25'b0000000000000100001101000;
    rom[197] = 25'b0000000000000100010100011;
    rom[198] = 25'b0000000000000100011011111;
    rom[199] = 25'b0000000000000100100011010;
    rom[200] = 25'b0000000000000100101010110;
    rom[201] = 25'b0000000000000100110010000;
    rom[202] = 25'b0000000000000100111001011;
    rom[203] = 25'b0000000000000101000000110;
    rom[204] = 25'b0000000000000101001000000;
    rom[205] = 25'b0000000000000101001111011;
    rom[206] = 25'b0000000000000101010110101;
    rom[207] = 25'b0000000000000101011101111;
    rom[208] = 25'b0000000000000101100101000;
    rom[209] = 25'b0000000000000101101100010;
    rom[210] = 25'b0000000000000101110011010;
    rom[211] = 25'b0000000000000101111010011;
    rom[212] = 25'b0000000000000110000001100;
    rom[213] = 25'b0000000000000110001000100;
    rom[214] = 25'b0000000000000110001111011;
    rom[215] = 25'b0000000000000110010110001;
    rom[216] = 25'b0000000000000110011101000;
    rom[217] = 25'b0000000000000110100011110;
    rom[218] = 25'b0000000000000110101010011;
    rom[219] = 25'b0000000000000110110000111;
    rom[220] = 25'b0000000000000110110111100;
    rom[221] = 25'b0000000000000110111101111;
    rom[222] = 25'b0000000000000111000100010;
    rom[223] = 25'b0000000000000111001010100;
    rom[224] = 25'b0000000000000111010000101;
    rom[225] = 25'b0000000000000111010110101;
    rom[226] = 25'b0000000000000111011100101;
    rom[227] = 25'b0000000000000111100010100;
    rom[228] = 25'b0000000000000111101000010;
    rom[229] = 25'b0000000000000111101101111;
    rom[230] = 25'b0000000000000111110011011;
    rom[231] = 25'b0000000000000111111000110;
    rom[232] = 25'b0000000000000111111110001;
    rom[233] = 25'b0000000000001000000011010;
    rom[234] = 25'b0000000000001000001000010;
    rom[235] = 25'b0000000000001000001101010;
    rom[236] = 25'b0000000000001000010010000;
    rom[237] = 25'b0000000000001000010110101;
    rom[238] = 25'b0000000000001000011011001;
    rom[239] = 25'b0000000000001000011111100;
    rom[240] = 25'b0000000000001000100011101;
    rom[241] = 25'b0000000000001000100111101;
    rom[242] = 25'b0000000000001000101011100;
    rom[243] = 25'b0000000000001000101111010;
    rom[244] = 25'b0000000000001000110010111;
    rom[245] = 25'b0000000000001000110110010;
    rom[246] = 25'b0000000000001000111001011;
    rom[247] = 25'b0000000000001000111100100;
    rom[248] = 25'b0000000000001000111111011;
    rom[249] = 25'b0000000000001001000010001;
    rom[250] = 25'b0000000000001001000100101;
    rom[251] = 25'b0000000000001001000110111;
    rom[252] = 25'b0000000000001001001001000;
    rom[253] = 25'b0000000000001001001010111;
    rom[254] = 25'b0000000000001001001100110;
    rom[255] = 25'b0000000000001001001110010;
    rom[256] = 25'b0000000000001001001111101;
    rom[257] = 25'b0000000000001001010000110;
    rom[258] = 25'b0000000000001001010001101;
    rom[259] = 25'b0000000000001001010010011;
    rom[260] = 25'b0000000000001001010010111;
    rom[261] = 25'b0000000000001001010011010;
    rom[262] = 25'b0000000000001001010011010;
    rom[263] = 25'b0000000000001001010011001;
    rom[264] = 25'b0000000000001001010010110;
    rom[265] = 25'b0000000000001001010010010;
    rom[266] = 25'b0000000000001001010001011;
    rom[267] = 25'b0000000000001001010000010;
    rom[268] = 25'b0000000000001001001111000;
    rom[269] = 25'b0000000000001001001101100;
    rom[270] = 25'b0000000000001001001011101;
    rom[271] = 25'b0000000000001001001001110;
    rom[272] = 25'b0000000000001001000111100;
    rom[273] = 25'b0000000000001001000101000;
    rom[274] = 25'b0000000000001001000010010;
    rom[275] = 25'b0000000000001000111111010;
    rom[276] = 25'b0000000000001000111100001;
    rom[277] = 25'b0000000000001000111000100;
    rom[278] = 25'b0000000000001000110100111;
    rom[279] = 25'b0000000000001000110000111;
    rom[280] = 25'b0000000000001000101100101;
    rom[281] = 25'b0000000000001000101000001;
    rom[282] = 25'b0000000000001000100011011;
    rom[283] = 25'b0000000000001000011110100;
    rom[284] = 25'b0000000000001000011001001;
    rom[285] = 25'b0000000000001000010011101;
    rom[286] = 25'b0000000000001000001101111;
    rom[287] = 25'b0000000000001000000111110;
    rom[288] = 25'b0000000000001000000001100;
    rom[289] = 25'b0000000000000111111011000;
    rom[290] = 25'b0000000000000111110100001;
    rom[291] = 25'b0000000000000111101101000;
    rom[292] = 25'b0000000000000111100101110;
    rom[293] = 25'b0000000000000111011110000;
    rom[294] = 25'b0000000000000111010110001;
    rom[295] = 25'b0000000000000111001110000;
    rom[296] = 25'b0000000000000111000101101;
    rom[297] = 25'b0000000000000110111101000;
    rom[298] = 25'b0000000000000110110100000;
    rom[299] = 25'b0000000000000110101010110;
    rom[300] = 25'b0000000000000110100001010;
    rom[301] = 25'b0000000000000110010111101;
    rom[302] = 25'b0000000000000110001101101;
    rom[303] = 25'b0000000000000110000011011;
    rom[304] = 25'b0000000000000101111000110;
    rom[305] = 25'b0000000000000101101110001;
    rom[306] = 25'b0000000000000101100011000;
    rom[307] = 25'b0000000000000101010111110;
    rom[308] = 25'b0000000000000101001100010;
    rom[309] = 25'b0000000000000101000000011;
    rom[310] = 25'b0000000000000100110100011;
    rom[311] = 25'b0000000000000100101000001;
    rom[312] = 25'b0000000000000100011011101;
    rom[313] = 25'b0000000000000100001110111;
    rom[314] = 25'b0000000000000100000001110;
    rom[315] = 25'b0000000000000011110100100;
    rom[316] = 25'b0000000000000011100111000;
    rom[317] = 25'b0000000000000011011001011;
    rom[318] = 25'b0000000000000011001011011;
    rom[319] = 25'b0000000000000010111101001;
    rom[320] = 25'b0000000000000010101110110;
    rom[321] = 25'b0000000000000010100000001;
    rom[322] = 25'b0000000000000010010001010;
    rom[323] = 25'b0000000000000010000010001;
    rom[324] = 25'b0000000000000001110010111;
    rom[325] = 25'b0000000000000001100011011;
    rom[326] = 25'b0000000000000001010011101;
    rom[327] = 25'b0000000000000001000011110;
    rom[328] = 25'b0000000000000000110011101;
    rom[329] = 25'b0000000000000000100011010;
    rom[330] = 25'b0000000000000000010010110;
    rom[331] = 25'b0000000000000000000010001;
    rom[332] = 25'b1111111111111111110001010;
    rom[333] = 25'b1111111111111111100000010;
    rom[334] = 25'b1111111111111111001111000;
    rom[335] = 25'b1111111111111110111101101;
    rom[336] = 25'b1111111111111110101100000;
    rom[337] = 25'b1111111111111110011010010;
    rom[338] = 25'b1111111111111110001000011;
    rom[339] = 25'b1111111111111101110110011;
    rom[340] = 25'b1111111111111101100100001;
    rom[341] = 25'b1111111111111101010001110;
    rom[342] = 25'b1111111111111100111111011;
    rom[343] = 25'b1111111111111100101100110;
    rom[344] = 25'b1111111111111100011010001;
    rom[345] = 25'b1111111111111100000111010;
    rom[346] = 25'b1111111111111011110100011;
    rom[347] = 25'b1111111111111011100001010;
    rom[348] = 25'b1111111111111011001110001;
    rom[349] = 25'b1111111111111010111010111;
    rom[350] = 25'b1111111111111010100111101;
    rom[351] = 25'b1111111111111010010100001;
    rom[352] = 25'b1111111111111010000000101;
    rom[353] = 25'b1111111111111001101101000;
    rom[354] = 25'b1111111111111001011001100;
    rom[355] = 25'b1111111111111001000101110;
    rom[356] = 25'b1111111111111000110010000;
    rom[357] = 25'b1111111111111000011110010;
    rom[358] = 25'b1111111111111000001010100;
    rom[359] = 25'b1111111111110111110110101;
    rom[360] = 25'b1111111111110111100010111;
    rom[361] = 25'b1111111111110111001111000;
    rom[362] = 25'b1111111111110110111011001;
    rom[363] = 25'b1111111111110110100111010;
    rom[364] = 25'b1111111111110110010011011;
    rom[365] = 25'b1111111111110101111111100;
    rom[366] = 25'b1111111111110101101011110;
    rom[367] = 25'b1111111111110101010111111;
    rom[368] = 25'b1111111111110101000100010;
    rom[369] = 25'b1111111111110100110000100;
    rom[370] = 25'b1111111111110100011100111;
    rom[371] = 25'b1111111111110100001001010;
    rom[372] = 25'b1111111111110011110101110;
    rom[373] = 25'b1111111111110011100010011;
    rom[374] = 25'b1111111111110011001111000;
    rom[375] = 25'b1111111111110010111011110;
    rom[376] = 25'b1111111111110010101000101;
    rom[377] = 25'b1111111111110010010101101;
    rom[378] = 25'b1111111111110010000010101;
    rom[379] = 25'b1111111111110001101111111;
    rom[380] = 25'b1111111111110001011101010;
    rom[381] = 25'b1111111111110001001010110;
    rom[382] = 25'b1111111111110000111000011;
    rom[383] = 25'b1111111111110000100110001;
    rom[384] = 25'b1111111111110000010100001;
    rom[385] = 25'b1111111111110000000010010;
    rom[386] = 25'b1111111111101111110000101;
    rom[387] = 25'b1111111111101111011111010;
    rom[388] = 25'b1111111111101111001110000;
    rom[389] = 25'b1111111111101110111100111;
    rom[390] = 25'b1111111111101110101100000;
    rom[391] = 25'b1111111111101110011011100;
    rom[392] = 25'b1111111111101110001011001;
    rom[393] = 25'b1111111111101101111011000;
    rom[394] = 25'b1111111111101101101011001;
    rom[395] = 25'b1111111111101101011011101;
    rom[396] = 25'b1111111111101101001100010;
    rom[397] = 25'b1111111111101100111101010;
    rom[398] = 25'b1111111111101100101110100;
    rom[399] = 25'b1111111111101100100000000;
    rom[400] = 25'b1111111111101100010001111;
    rom[401] = 25'b1111111111101100000100001;
    rom[402] = 25'b1111111111101011110110101;
    rom[403] = 25'b1111111111101011101001011;
    rom[404] = 25'b1111111111101011011100100;
    rom[405] = 25'b1111111111101011010000001;
    rom[406] = 25'b1111111111101011000100000;
    rom[407] = 25'b1111111111101010111000010;
    rom[408] = 25'b1111111111101010101100111;
    rom[409] = 25'b1111111111101010100001110;
    rom[410] = 25'b1111111111101010010111001;
    rom[411] = 25'b1111111111101010001101000;
    rom[412] = 25'b1111111111101010000011001;
    rom[413] = 25'b1111111111101001111001101;
    rom[414] = 25'b1111111111101001110000110;
    rom[415] = 25'b1111111111101001101000001;
    rom[416] = 25'b1111111111101001100000000;
    rom[417] = 25'b1111111111101001011000010;
    rom[418] = 25'b1111111111101001010001001;
    rom[419] = 25'b1111111111101001001010010;
    rom[420] = 25'b1111111111101001000100000;
    rom[421] = 25'b1111111111101000111110001;
    rom[422] = 25'b1111111111101000111000110;
    rom[423] = 25'b1111111111101000110011111;
    rom[424] = 25'b1111111111101000101111100;
    rom[425] = 25'b1111111111101000101011100;
    rom[426] = 25'b1111111111101000101000010;
    rom[427] = 25'b1111111111101000100101010;
    rom[428] = 25'b1111111111101000100011000;
    rom[429] = 25'b1111111111101000100001001;
    rom[430] = 25'b1111111111101000011111110;
    rom[431] = 25'b1111111111101000011111000;
    rom[432] = 25'b1111111111101000011110110;
    rom[433] = 25'b1111111111101000011111000;
    rom[434] = 25'b1111111111101000011111111;
    rom[435] = 25'b1111111111101000100001010;
    rom[436] = 25'b1111111111101000100011011;
    rom[437] = 25'b1111111111101000100101111;
    rom[438] = 25'b1111111111101000101000111;
    rom[439] = 25'b1111111111101000101100101;
    rom[440] = 25'b1111111111101000110001000;
    rom[441] = 25'b1111111111101000110101110;
    rom[442] = 25'b1111111111101000111011010;
    rom[443] = 25'b1111111111101001000001010;
    rom[444] = 25'b1111111111101001000111111;
    rom[445] = 25'b1111111111101001001111000;
    rom[446] = 25'b1111111111101001010110111;
    rom[447] = 25'b1111111111101001011111011;
    rom[448] = 25'b1111111111101001101000011;
    rom[449] = 25'b1111111111101001110010001;
    rom[450] = 25'b1111111111101001111100011;
    rom[451] = 25'b1111111111101010000111010;
    rom[452] = 25'b1111111111101010010010110;
    rom[453] = 25'b1111111111101010011110111;
    rom[454] = 25'b1111111111101010101011101;
    rom[455] = 25'b1111111111101010111001000;
    rom[456] = 25'b1111111111101011000111000;
    rom[457] = 25'b1111111111101011010101101;
    rom[458] = 25'b1111111111101011100100111;
    rom[459] = 25'b1111111111101011110100110;
    rom[460] = 25'b1111111111101100000101010;
    rom[461] = 25'b1111111111101100010110011;
    rom[462] = 25'b1111111111101100101000001;
    rom[463] = 25'b1111111111101100111010100;
    rom[464] = 25'b1111111111101101001101100;
    rom[465] = 25'b1111111111101101100001010;
    rom[466] = 25'b1111111111101101110101011;
    rom[467] = 25'b1111111111101110001010011;
    rom[468] = 25'b1111111111101110011111111;
    rom[469] = 25'b1111111111101110110110000;
    rom[470] = 25'b1111111111101111001100110;
    rom[471] = 25'b1111111111101111100100001;
    rom[472] = 25'b1111111111101111111100001;
    rom[473] = 25'b1111111111110000010100101;
    rom[474] = 25'b1111111111110000101101111;
    rom[475] = 25'b1111111111110001000111110;
    rom[476] = 25'b1111111111110001100010001;
    rom[477] = 25'b1111111111110001111101000;
    rom[478] = 25'b1111111111110010011000101;
    rom[479] = 25'b1111111111110010110100111;
    rom[480] = 25'b1111111111110011010001101;
    rom[481] = 25'b1111111111110011101111000;
    rom[482] = 25'b1111111111110100001100111;
    rom[483] = 25'b1111111111110100101011011;
    rom[484] = 25'b1111111111110101001010011;
    rom[485] = 25'b1111111111110101101010000;
    rom[486] = 25'b1111111111110110001010001;
    rom[487] = 25'b1111111111110110101010111;
    rom[488] = 25'b1111111111110111001100001;
    rom[489] = 25'b1111111111110111101101111;
    rom[490] = 25'b1111111111111000010000010;
    rom[491] = 25'b1111111111111000110011000;
    rom[492] = 25'b1111111111111001010110010;
    rom[493] = 25'b1111111111111001111010001;
    rom[494] = 25'b1111111111111010011110100;
    rom[495] = 25'b1111111111111011000011010;
    rom[496] = 25'b1111111111111011101000100;
    rom[497] = 25'b1111111111111100001110010;
    rom[498] = 25'b1111111111111100110100011;
    rom[499] = 25'b1111111111111101011011000;
    rom[500] = 25'b1111111111111110000010001;
    rom[501] = 25'b1111111111111110101001100;
    rom[502] = 25'b1111111111111111010001011;
    rom[503] = 25'b1111111111111111111001110;
    rom[504] = 25'b0000000000000000100010011;
    rom[505] = 25'b0000000000000001001011100;
    rom[506] = 25'b0000000000000001110100111;
    rom[507] = 25'b0000000000000010011110110;
    rom[508] = 25'b0000000000000011001000111;
    rom[509] = 25'b0000000000000011110011011;
    rom[510] = 25'b0000000000000100011110010;
    rom[511] = 25'b0000000000000101001001011;
    rom[512] = 25'b0000000000000101110100110;
    rom[513] = 25'b0000000000000110100000101;
    rom[514] = 25'b0000000000000111001100101;
    rom[515] = 25'b0000000000000111111000110;
    rom[516] = 25'b0000000000001000100101011;
    rom[517] = 25'b0000000000001001010010001;
    rom[518] = 25'b0000000000001001111111000;
    rom[519] = 25'b0000000000001010101100001;
    rom[520] = 25'b0000000000001011011001100;
    rom[521] = 25'b0000000000001100000111000;
    rom[522] = 25'b0000000000001100110100110;
    rom[523] = 25'b0000000000001101100010100;
    rom[524] = 25'b0000000000001110010000011;
    rom[525] = 25'b0000000000001110111110100;
    rom[526] = 25'b0000000000001111101100101;
    rom[527] = 25'b0000000000010000011010111;
    rom[528] = 25'b0000000000010001001001001;
    rom[529] = 25'b0000000000010001110111011;
    rom[530] = 25'b0000000000010010100101111;
    rom[531] = 25'b0000000000010011010100001;
    rom[532] = 25'b0000000000010100000010101;
    rom[533] = 25'b0000000000010100110000111;
    rom[534] = 25'b0000000000010101011111010;
    rom[535] = 25'b0000000000010110001101100;
    rom[536] = 25'b0000000000010110111011110;
    rom[537] = 25'b0000000000010111101001111;
    rom[538] = 25'b0000000000011000010111111;
    rom[539] = 25'b0000000000011001000101101;
    rom[540] = 25'b0000000000011001110011100;
    rom[541] = 25'b0000000000011010100001000;
    rom[542] = 25'b0000000000011011001110011;
    rom[543] = 25'b0000000000011011111011100;
    rom[544] = 25'b0000000000011100101000101;
    rom[545] = 25'b0000000000011101010101011;
    rom[546] = 25'b0000000000011110000001110;
    rom[547] = 25'b0000000000011110101110000;
    rom[548] = 25'b0000000000011111011010000;
    rom[549] = 25'b0000000000100000000101101;
    rom[550] = 25'b0000000000100000110000111;
    rom[551] = 25'b0000000000100001011011110;
    rom[552] = 25'b0000000000100010000110011;
    rom[553] = 25'b0000000000100010110000100;
    rom[554] = 25'b0000000000100011011010011;
    rom[555] = 25'b0000000000100100000011110;
    rom[556] = 25'b0000000000100100101100110;
    rom[557] = 25'b0000000000100101010101001;
    rom[558] = 25'b0000000000100101111101001;
    rom[559] = 25'b0000000000100110100100101;
    rom[560] = 25'b0000000000100111001011100;
    rom[561] = 25'b0000000000100111110010000;
    rom[562] = 25'b0000000000101000010111111;
    rom[563] = 25'b0000000000101000111101001;
    rom[564] = 25'b0000000000101001100001111;
    rom[565] = 25'b0000000000101010000110000;
    rom[566] = 25'b0000000000101010101001011;
    rom[567] = 25'b0000000000101011001100010;
    rom[568] = 25'b0000000000101011101110011;
    rom[569] = 25'b0000000000101100001111111;
    rom[570] = 25'b0000000000101100110000101;
    rom[571] = 25'b0000000000101101010000100;
    rom[572] = 25'b0000000000101101101111111;
    rom[573] = 25'b0000000000101110001110011;
    rom[574] = 25'b0000000000101110101100001;
    rom[575] = 25'b0000000000101111001001000;
    rom[576] = 25'b0000000000101111100101001;
    rom[577] = 25'b0000000000110000000000100;
    rom[578] = 25'b0000000000110000011010111;
    rom[579] = 25'b0000000000110000110100011;
    rom[580] = 25'b0000000000110001001101001;
    rom[581] = 25'b0000000000110001100100111;
    rom[582] = 25'b0000000000110001111011101;
    rom[583] = 25'b0000000000110010010001101;
    rom[584] = 25'b0000000000110010100110100;
    rom[585] = 25'b0000000000110010111010100;
    rom[586] = 25'b0000000000110011001101011;
    rom[587] = 25'b0000000000110011011111011;
    rom[588] = 25'b0000000000110011110000011;
    rom[589] = 25'b0000000000110100000000011;
    rom[590] = 25'b0000000000110100001111010;
    rom[591] = 25'b0000000000110100011101000;
    rom[592] = 25'b0000000000110100101001110;
    rom[593] = 25'b0000000000110100110101011;
    rom[594] = 25'b0000000000110100111111111;
    rom[595] = 25'b0000000000110101001001010;
    rom[596] = 25'b0000000000110101010001100;
    rom[597] = 25'b0000000000110101011000110;
    rom[598] = 25'b0000000000110101011110100;
    rom[599] = 25'b0000000000110101100011011;
    rom[600] = 25'b0000000000110101100111000;
    rom[601] = 25'b0000000000110101101001011;
    rom[602] = 25'b0000000000110101101010100;
    rom[603] = 25'b0000000000110101101010011;
    rom[604] = 25'b0000000000110101101001001;
    rom[605] = 25'b0000000000110101100110101;
    rom[606] = 25'b0000000000110101100010110;
    rom[607] = 25'b0000000000110101011101110;
    rom[608] = 25'b0000000000110101010111011;
    rom[609] = 25'b0000000000110101001111110;
    rom[610] = 25'b0000000000110101000110110;
    rom[611] = 25'b0000000000110100111100100;
    rom[612] = 25'b0000000000110100110001000;
    rom[613] = 25'b0000000000110100100100001;
    rom[614] = 25'b0000000000110100010110000;
    rom[615] = 25'b0000000000110100000110011;
    rom[616] = 25'b0000000000110011110101100;
    rom[617] = 25'b0000000000110011100011010;
    rom[618] = 25'b0000000000110011001111101;
    rom[619] = 25'b0000000000110010111010110;
    rom[620] = 25'b0000000000110010100100011;
    rom[621] = 25'b0000000000110010001100110;
    rom[622] = 25'b0000000000110001110011110;
    rom[623] = 25'b0000000000110001011001010;
    rom[624] = 25'b0000000000110000111101100;
    rom[625] = 25'b0000000000110000100000011;
    rom[626] = 25'b0000000000110000000001110;
    rom[627] = 25'b0000000000101111100001111;
    rom[628] = 25'b0000000000101111000000100;
    rom[629] = 25'b0000000000101110011101111;
    rom[630] = 25'b0000000000101101111001110;
    rom[631] = 25'b0000000000101101010100001;
    rom[632] = 25'b0000000000101100101101011;
    rom[633] = 25'b0000000000101100000101001;
    rom[634] = 25'b0000000000101011011011100;
    rom[635] = 25'b0000000000101010110000100;
    rom[636] = 25'b0000000000101010000100001;
    rom[637] = 25'b0000000000101001010110011;
    rom[638] = 25'b0000000000101000100111010;
    rom[639] = 25'b0000000000100111110110110;
    rom[640] = 25'b0000000000100111000100111;
    rom[641] = 25'b0000000000100110010001110;
    rom[642] = 25'b0000000000100101011101010;
    rom[643] = 25'b0000000000100100100111011;
    rom[644] = 25'b0000000000100011110000010;
    rom[645] = 25'b0000000000100010110111110;
    rom[646] = 25'b0000000000100001111101111;
    rom[647] = 25'b0000000000100001000010111;
    rom[648] = 25'b0000000000100000000110011;
    rom[649] = 25'b0000000000011111001000110;
    rom[650] = 25'b0000000000011110001001110;
    rom[651] = 25'b0000000000011101001001101;
    rom[652] = 25'b0000000000011100001000000;
    rom[653] = 25'b0000000000011011000101011;
    rom[654] = 25'b0000000000011010000001011;
    rom[655] = 25'b0000000000011000111100010;
    rom[656] = 25'b0000000000010111110110000;
    rom[657] = 25'b0000000000010110101110100;
    rom[658] = 25'b0000000000010101100101110;
    rom[659] = 25'b0000000000010100011100000;
    rom[660] = 25'b0000000000010011010001000;
    rom[661] = 25'b0000000000010010000101000;
    rom[662] = 25'b0000000000010000110111110;
    rom[663] = 25'b0000000000001111101001100;
    rom[664] = 25'b0000000000001110011010010;
    rom[665] = 25'b0000000000001101001001111;
    rom[666] = 25'b0000000000001011111000100;
    rom[667] = 25'b0000000000001010100110001;
    rom[668] = 25'b0000000000001001010010111;
    rom[669] = 25'b0000000000000111111110100;
    rom[670] = 25'b0000000000000110101001010;
    rom[671] = 25'b0000000000000101010011001;
    rom[672] = 25'b0000000000000011111100001;
    rom[673] = 25'b0000000000000010100100001;
    rom[674] = 25'b0000000000000001001011100;
    rom[675] = 25'b1111111111111111110010000;
    rom[676] = 25'b1111111111111110010111101;
    rom[677] = 25'b1111111111111100111100100;
    rom[678] = 25'b1111111111111011100000101;
    rom[679] = 25'b1111111111111010000100000;
    rom[680] = 25'b1111111111111000100110110;
    rom[681] = 25'b1111111111110111001000110;
    rom[682] = 25'b1111111111110101101010010;
    rom[683] = 25'b1111111111110100001011001;
    rom[684] = 25'b1111111111110010101011011;
    rom[685] = 25'b1111111111110001001011001;
    rom[686] = 25'b1111111111101111101010011;
    rom[687] = 25'b1111111111101110001001001;
    rom[688] = 25'b1111111111101100100111011;
    rom[689] = 25'b1111111111101011000101010;
    rom[690] = 25'b1111111111101001100010110;
    rom[691] = 25'b1111111111100111111111111;
    rom[692] = 25'b1111111111100110011100101;
    rom[693] = 25'b1111111111100100111001001;
    rom[694] = 25'b1111111111100011010101100;
    rom[695] = 25'b1111111111100001110001011;
    rom[696] = 25'b1111111111100000001101010;
    rom[697] = 25'b1111111111011110101000111;
    rom[698] = 25'b1111111111011101000100100;
    rom[699] = 25'b1111111111011011100000000;
    rom[700] = 25'b1111111111011001111011100;
    rom[701] = 25'b1111111111011000010110111;
    rom[702] = 25'b1111111111010110110010010;
    rom[703] = 25'b1111111111010101001101110;
    rom[704] = 25'b1111111111010011101001011;
    rom[705] = 25'b1111111111010010000101010;
    rom[706] = 25'b1111111111010000100001001;
    rom[707] = 25'b1111111111001110111101010;
    rom[708] = 25'b1111111111001101011001101;
    rom[709] = 25'b1111111111001011110110010;
    rom[710] = 25'b1111111111001010010011010;
    rom[711] = 25'b1111111111001000110000100;
    rom[712] = 25'b1111111111000111001110010;
    rom[713] = 25'b1111111111000101101100100;
    rom[714] = 25'b1111111111000100001011001;
    rom[715] = 25'b1111111111000010101010011;
    rom[716] = 25'b1111111111000001001010001;
    rom[717] = 25'b1111111110111111101010100;
    rom[718] = 25'b1111111110111110001011011;
    rom[719] = 25'b1111111110111100101101000;
    rom[720] = 25'b1111111110111011001111100;
    rom[721] = 25'b1111111110111001110010101;
    rom[722] = 25'b1111111110111000010110100;
    rom[723] = 25'b1111111110110110111011011;
    rom[724] = 25'b1111111110110101100001000;
    rom[725] = 25'b1111111110110100000111100;
    rom[726] = 25'b1111111110110010101111001;
    rom[727] = 25'b1111111110110001010111101;
    rom[728] = 25'b1111111110110000000001001;
    rom[729] = 25'b1111111110101110101011111;
    rom[730] = 25'b1111111110101101010111101;
    rom[731] = 25'b1111111110101100000100100;
    rom[732] = 25'b1111111110101010110010101;
    rom[733] = 25'b1111111110101001100010000;
    rom[734] = 25'b1111111110101000010010101;
    rom[735] = 25'b1111111110100111000100101;
    rom[736] = 25'b1111111110100101111000000;
    rom[737] = 25'b1111111110100100101100101;
    rom[738] = 25'b1111111110100011100010111;
    rom[739] = 25'b1111111110100010011010100;
    rom[740] = 25'b1111111110100001010011101;
    rom[741] = 25'b1111111110100000001110010;
    rom[742] = 25'b1111111110011111001010101;
    rom[743] = 25'b1111111110011110001000100;
    rom[744] = 25'b1111111110011101001000001;
    rom[745] = 25'b1111111110011100001001100;
    rom[746] = 25'b1111111110011011001100100;
    rom[747] = 25'b1111111110011010010001011;
    rom[748] = 25'b1111111110011001010111111;
    rom[749] = 25'b1111111110011000100000100;
    rom[750] = 25'b1111111110010111101010110;
    rom[751] = 25'b1111111110010110110111001;
    rom[752] = 25'b1111111110010110000101011;
    rom[753] = 25'b1111111110010101010101101;
    rom[754] = 25'b1111111110010100100111111;
    rom[755] = 25'b1111111110010011111100010;
    rom[756] = 25'b1111111110010011010010101;
    rom[757] = 25'b1111111110010010101011010;
    rom[758] = 25'b1111111110010010000101111;
    rom[759] = 25'b1111111110010001100010110;
    rom[760] = 25'b1111111110010001000001111;
    rom[761] = 25'b1111111110010000100011010;
    rom[762] = 25'b1111111110010000000111000;
    rom[763] = 25'b1111111110001111101100111;
    rom[764] = 25'b1111111110001111010101001;
    rom[765] = 25'b1111111110001110111111111;
    rom[766] = 25'b1111111110001110101101000;
    rom[767] = 25'b1111111110001110011100100;
    rom[768] = 25'b1111111110001110001110011;
    rom[769] = 25'b1111111110001110000010111;
    rom[770] = 25'b1111111110001101111001110;
    rom[771] = 25'b1111111110001101110011010;
    rom[772] = 25'b1111111110001101101111010;
    rom[773] = 25'b1111111110001101101101110;
    rom[774] = 25'b1111111110001101101111000;
    rom[775] = 25'b1111111110001101110010110;
    rom[776] = 25'b1111111110001101111001001;
    rom[777] = 25'b1111111110001110000010011;
    rom[778] = 25'b1111111110001110001110000;
    rom[779] = 25'b1111111110001110011100100;
    rom[780] = 25'b1111111110001110101101101;
    rom[781] = 25'b1111111110001111000001100;
    rom[782] = 25'b1111111110001111011000001;
    rom[783] = 25'b1111111110001111110001100;
    rom[784] = 25'b1111111110010000001101110;
    rom[785] = 25'b1111111110010000101100110;
    rom[786] = 25'b1111111110010001001110100;
    rom[787] = 25'b1111111110010001110011000;
    rom[788] = 25'b1111111110010010011010011;
    rom[789] = 25'b1111111110010011000100101;
    rom[790] = 25'b1111111110010011110001101;
    rom[791] = 25'b1111111110010100100001100;
    rom[792] = 25'b1111111110010101010100010;
    rom[793] = 25'b1111111110010110001001110;
    rom[794] = 25'b1111111110010111000010010;
    rom[795] = 25'b1111111110010111111101101;
    rom[796] = 25'b1111111110011000111011110;
    rom[797] = 25'b1111111110011001111100111;
    rom[798] = 25'b1111111110011011000000110;
    rom[799] = 25'b1111111110011100000111100;
    rom[800] = 25'b1111111110011101010001001;
    rom[801] = 25'b1111111110011110011101110;
    rom[802] = 25'b1111111110011111101101001;
    rom[803] = 25'b1111111110100000111111011;
    rom[804] = 25'b1111111110100010010100100;
    rom[805] = 25'b1111111110100011101100011;
    rom[806] = 25'b1111111110100101000111001;
    rom[807] = 25'b1111111110100110100100110;
    rom[808] = 25'b1111111110101000000101001;
    rom[809] = 25'b1111111110101001101000010;
    rom[810] = 25'b1111111110101011001110011;
    rom[811] = 25'b1111111110101100110111001;
    rom[812] = 25'b1111111110101110100010110;
    rom[813] = 25'b1111111110110000010001000;
    rom[814] = 25'b1111111110110010000010000;
    rom[815] = 25'b1111111110110011110101110;
    rom[816] = 25'b1111111110110101101100010;
    rom[817] = 25'b1111111110110111100101011;
    rom[818] = 25'b1111111110111001100001001;
    rom[819] = 25'b1111111110111011011111011;
    rom[820] = 25'b1111111110111101100000011;
    rom[821] = 25'b1111111110111111100100000;
    rom[822] = 25'b1111111111000001101010001;
    rom[823] = 25'b1111111111000011110010111;
    rom[824] = 25'b1111111111000101111110000;
    rom[825] = 25'b1111111111001000001011101;
    rom[826] = 25'b1111111111001010011011101;
    rom[827] = 25'b1111111111001100101110001;
    rom[828] = 25'b1111111111001111000011000;
    rom[829] = 25'b1111111111010001011010010;
    rom[830] = 25'b1111111111010011110011101;
    rom[831] = 25'b1111111111010110001111011;
    rom[832] = 25'b1111111111011000101101011;
    rom[833] = 25'b1111111111011011001101101;
    rom[834] = 25'b1111111111011101110000000;
    rom[835] = 25'b1111111111100000010100011;
    rom[836] = 25'b1111111111100010111011000;
    rom[837] = 25'b1111111111100101100011100;
    rom[838] = 25'b1111111111101000001110001;
    rom[839] = 25'b1111111111101010111010100;
    rom[840] = 25'b1111111111101101101001000;
    rom[841] = 25'b1111111111110000011001001;
    rom[842] = 25'b1111111111110011001011001;
    rom[843] = 25'b1111111111110101111111000;
    rom[844] = 25'b1111111111111000110100011;
    rom[845] = 25'b1111111111111011101011100;
    rom[846] = 25'b1111111111111110100100010;
    rom[847] = 25'b0000000000000001011110100;
    rom[848] = 25'b0000000000000100011010010;
    rom[849] = 25'b0000000000000111010111011;
    rom[850] = 25'b0000000000001010010101111;
    rom[851] = 25'b0000000000001101010101110;
    rom[852] = 25'b0000000000010000010111000;
    rom[853] = 25'b0000000000010011011001010;
    rom[854] = 25'b0000000000010110011100110;
    rom[855] = 25'b0000000000011001100001010;
    rom[856] = 25'b0000000000011100100110111;
    rom[857] = 25'b0000000000011111101101100;
    rom[858] = 25'b0000000000100010110100111;
    rom[859] = 25'b0000000000100101111101001;
    rom[860] = 25'b0000000000101001000110001;
    rom[861] = 25'b0000000000101100001111111;
    rom[862] = 25'b0000000000101111011010010;
    rom[863] = 25'b0000000000110010100101001;
    rom[864] = 25'b0000000000110101110000100;
    rom[865] = 25'b0000000000111000111100011;
    rom[866] = 25'b0000000000111100001000101;
    rom[867] = 25'b0000000000111111010101001;
    rom[868] = 25'b0000000001000010100001110;
    rom[869] = 25'b0000000001000101101110101;
    rom[870] = 25'b0000000001001000111011100;
    rom[871] = 25'b0000000001001100001000100;
    rom[872] = 25'b0000000001001111010101011;
    rom[873] = 25'b0000000001010010100010001;
    rom[874] = 25'b0000000001010101101110100;
    rom[875] = 25'b0000000001011000111010110;
    rom[876] = 25'b0000000001011100000110101;
    rom[877] = 25'b0000000001011111010010000;
    rom[878] = 25'b0000000001100010011100110;
    rom[879] = 25'b0000000001100101100111001;
    rom[880] = 25'b0000000001101000110000101;
    rom[881] = 25'b0000000001101011111001011;
    rom[882] = 25'b0000000001101111000001011;
    rom[883] = 25'b0000000001110010001000100;
    rom[884] = 25'b0000000001110101001110100;
    rom[885] = 25'b0000000001111000010011100;
    rom[886] = 25'b0000000001111011010111011;
    rom[887] = 25'b0000000001111110011010000;
    rom[888] = 25'b0000000010000001011011011;
    rom[889] = 25'b0000000010000100011011010;
    rom[890] = 25'b0000000010000111011001110;
    rom[891] = 25'b0000000010001010010110101;
    rom[892] = 25'b0000000010001101010001111;
    rom[893] = 25'b0000000010010000001011100;
    rom[894] = 25'b0000000010010011000011011;
    rom[895] = 25'b0000000010010101111001010;
    rom[896] = 25'b0000000010011000101101010;
    rom[897] = 25'b0000000010011011011111010;
    rom[898] = 25'b0000000010011110001111000;
    rom[899] = 25'b0000000010100000111100110;
    rom[900] = 25'b0000000010100011101000001;
    rom[901] = 25'b0000000010100110010001010;
    rom[902] = 25'b0000000010101000110111111;
    rom[903] = 25'b0000000010101011011100000;
    rom[904] = 25'b0000000010101101111101101;
    rom[905] = 25'b0000000010110000011100100;
    rom[906] = 25'b0000000010110010111000101;
    rom[907] = 25'b0000000010110101010010000;
    rom[908] = 25'b0000000010110111101000100;
    rom[909] = 25'b0000000010111001111100000;
    rom[910] = 25'b0000000010111100001100011;
    rom[911] = 25'b0000000010111110011001111;
    rom[912] = 25'b0000000011000000100100000;
    rom[913] = 25'b0000000011000010101010111;
    rom[914] = 25'b0000000011000100101110011;
    rom[915] = 25'b0000000011000110101110100;
    rom[916] = 25'b0000000011001000101011001;
    rom[917] = 25'b0000000011001010100100010;
    rom[918] = 25'b0000000011001100011001101;
    rom[919] = 25'b0000000011001110001011011;
    rom[920] = 25'b0000000011001111111001011;
    rom[921] = 25'b0000000011010001100011100;
    rom[922] = 25'b0000000011010011001001110;
    rom[923] = 25'b0000000011010100101100000;
    rom[924] = 25'b0000000011010110001010010;
    rom[925] = 25'b0000000011010111100100011;
    rom[926] = 25'b0000000011011000111010010;
    rom[927] = 25'b0000000011011010001100000;
    rom[928] = 25'b0000000011011011011001011;
    rom[929] = 25'b0000000011011100100010100;
    rom[930] = 25'b0000000011011101100111001;
    rom[931] = 25'b0000000011011110100111010;
    rom[932] = 25'b0000000011011111100010111;
    rom[933] = 25'b0000000011100000011001111;
    rom[934] = 25'b0000000011100001001100010;
    rom[935] = 25'b0000000011100001111010000;
    rom[936] = 25'b0000000011100010100010111;
    rom[937] = 25'b0000000011100011000111001;
    rom[938] = 25'b0000000011100011100110011;
    rom[939] = 25'b0000000011100100000000110;
    rom[940] = 25'b0000000011100100010110010;
    rom[941] = 25'b0000000011100100100110101;
    rom[942] = 25'b0000000011100100110010000;
    rom[943] = 25'b0000000011100100111000011;
    rom[944] = 25'b0000000011100100111001100;
    rom[945] = 25'b0000000011100100110101100;
    rom[946] = 25'b0000000011100100101100010;
    rom[947] = 25'b0000000011100100011101111;
    rom[948] = 25'b0000000011100100001010001;
    rom[949] = 25'b0000000011100011110001001;
    rom[950] = 25'b0000000011100011010010111;
    rom[951] = 25'b0000000011100010101111000;
    rom[952] = 25'b0000000011100010000101111;
    rom[953] = 25'b0000000011100001010111010;
    rom[954] = 25'b0000000011100000100011010;
    rom[955] = 25'b0000000011011111101001110;
    rom[956] = 25'b0000000011011110101010110;
    rom[957] = 25'b0000000011011101100110010;
    rom[958] = 25'b0000000011011100011100010;
    rom[959] = 25'b0000000011011011001100101;
    rom[960] = 25'b0000000011011001110111011;
    rom[961] = 25'b0000000011011000011100101;
    rom[962] = 25'b0000000011010110111100011;
    rom[963] = 25'b0000000011010101010110011;
    rom[964] = 25'b0000000011010011101010110;
    rom[965] = 25'b0000000011010001111001101;
    rom[966] = 25'b0000000011010000000010111;
    rom[967] = 25'b0000000011001110000110011;
    rom[968] = 25'b0000000011001100000100100;
    rom[969] = 25'b0000000011001001111100111;
    rom[970] = 25'b0000000011000111101111101;
    rom[971] = 25'b0000000011000101011100111;
    rom[972] = 25'b0000000011000011000100010;
    rom[973] = 25'b0000000011000000100110011;
    rom[974] = 25'b0000000010111110000010110;
    rom[975] = 25'b0000000010111011011001110;
    rom[976] = 25'b0000000010111000101011001;
    rom[977] = 25'b0000000010110101110110111;
    rom[978] = 25'b0000000010110010111101011;
    rom[979] = 25'b0000000010101111111110010;
    rom[980] = 25'b0000000010101100111001110;
    rom[981] = 25'b0000000010101001101111111;
    rom[982] = 25'b0000000010100110100000100;
    rom[983] = 25'b0000000010100011001011111;
    rom[984] = 25'b0000000010011111110010000;
    rom[985] = 25'b0000000010011100010010110;
    rom[986] = 25'b0000000010011000101110010;
    rom[987] = 25'b0000000010010101000100101;
    rom[988] = 25'b0000000010010001010101110;
    rom[989] = 25'b0000000010001101100001111;
    rom[990] = 25'b0000000010001001101001000;
    rom[991] = 25'b0000000010000101101011000;
    rom[992] = 25'b0000000010000001101000001;
    rom[993] = 25'b0000000001111101100000010;
    rom[994] = 25'b0000000001111001010011101;
    rom[995] = 25'b0000000001110101000010010;
    rom[996] = 25'b0000000001110000101100001;
    rom[997] = 25'b0000000001101100010001011;
    rom[998] = 25'b0000000001100111110010000;
    rom[999] = 25'b0000000001100011001110001;
    rom[1000] = 25'b0000000001011110100101110;
    rom[1001] = 25'b0000000001011001111001001;
    rom[1002] = 25'b0000000001010101001000000;
    rom[1003] = 25'b0000000001010000010010101;
    rom[1004] = 25'b0000000001001011011001010;
    rom[1005] = 25'b0000000001000110011011110;
    rom[1006] = 25'b0000000001000001011010011;
    rom[1007] = 25'b0000000000111100010101000;
    rom[1008] = 25'b0000000000110111001011110;
    rom[1009] = 25'b0000000000110001111110111;
    rom[1010] = 25'b0000000000101100101110010;
    rom[1011] = 25'b0000000000100111011010001;
    rom[1012] = 25'b0000000000100010000010100;
    rom[1013] = 25'b0000000000011100100111101;
    rom[1014] = 25'b0000000000010111001001011;
    rom[1015] = 25'b0000000000010001101000000;
    rom[1016] = 25'b0000000000001100000011101;
    rom[1017] = 25'b0000000000000110011100010;
    rom[1018] = 25'b0000000000000000110010001;
    rom[1019] = 25'b1111111111111011000101010;
    rom[1020] = 25'b1111111111110101010101101;
    rom[1021] = 25'b1111111111101111100011100;
    rom[1022] = 25'b1111111111101001101111000;
    rom[1023] = 25'b1111111111100011111000010;
    rom[1024] = 25'b1111111111011101111111001;
    rom[1025] = 25'b1111111111011000000100001;
    rom[1026] = 25'b1111111111010010000111001;
    rom[1027] = 25'b1111111111001100001000011;
    rom[1028] = 25'b1111111111000110000111110;
    rom[1029] = 25'b1111111111000000000101110;
    rom[1030] = 25'b1111111110111010000010010;
    rom[1031] = 25'b1111111110110011111101011;
    rom[1032] = 25'b1111111110101101110111010;
    rom[1033] = 25'b1111111110100111110000010;
    rom[1034] = 25'b1111111110100001101000001;
    rom[1035] = 25'b1111111110011011011111011;
    rom[1036] = 25'b1111111110010101010101110;
    rom[1037] = 25'b1111111110001111001011110;
    rom[1038] = 25'b1111111110001001000001010;
    rom[1039] = 25'b1111111110000010110110101;
    rom[1040] = 25'b1111111101111100101011111;
    rom[1041] = 25'b1111111101110110100001000;
    rom[1042] = 25'b1111111101110000010110011;
    rom[1043] = 25'b1111111101101010001100000;
    rom[1044] = 25'b1111111101100100000010001;
    rom[1045] = 25'b1111111101011101111000110;
    rom[1046] = 25'b1111111101010111110000010;
    rom[1047] = 25'b1111111101010001101000100;
    rom[1048] = 25'b1111111101001011100001110;
    rom[1049] = 25'b1111111101000101011100010;
    rom[1050] = 25'b1111111100111111011000000;
    rom[1051] = 25'b1111111100111001010101010;
    rom[1052] = 25'b1111111100110011010100000;
    rom[1053] = 25'b1111111100101101010100101;
    rom[1054] = 25'b1111111100100111010111010;
    rom[1055] = 25'b1111111100100001011011110;
    rom[1056] = 25'b1111111100011011100010100;
    rom[1057] = 25'b1111111100010101101011101;
    rom[1058] = 25'b1111111100001111110111001;
    rom[1059] = 25'b1111111100001010000101100;
    rom[1060] = 25'b1111111100000100010110101;
    rom[1061] = 25'b1111111011111110101010101;
    rom[1062] = 25'b1111111011111001000001110;
    rom[1063] = 25'b1111111011110011011100000;
    rom[1064] = 25'b1111111011101101111001111;
    rom[1065] = 25'b1111111011101000011011010;
    rom[1066] = 25'b1111111011100011000000010;
    rom[1067] = 25'b1111111011011101101001001;
    rom[1068] = 25'b1111111011011000010110001;
    rom[1069] = 25'b1111111011010011000111010;
    rom[1070] = 25'b1111111011001101111100101;
    rom[1071] = 25'b1111111011001000110110011;
    rom[1072] = 25'b1111111011000011110100110;
    rom[1073] = 25'b1111111010111110111000000;
    rom[1074] = 25'b1111111010111010000000001;
    rom[1075] = 25'b1111111010110101001101010;
    rom[1076] = 25'b1111111010110000011111100;
    rom[1077] = 25'b1111111010101011110111001;
    rom[1078] = 25'b1111111010100111010100010;
    rom[1079] = 25'b1111111010100010110111000;
    rom[1080] = 25'b1111111010011110011111100;
    rom[1081] = 25'b1111111010011010001101111;
    rom[1082] = 25'b1111111010010110000010011;
    rom[1083] = 25'b1111111010010001111101000;
    rom[1084] = 25'b1111111010001101111110000;
    rom[1085] = 25'b1111111010001010000101011;
    rom[1086] = 25'b1111111010000110010011011;
    rom[1087] = 25'b1111111010000010101000001;
    rom[1088] = 25'b1111111001111111000011101;
    rom[1089] = 25'b1111111001111011100110001;
    rom[1090] = 25'b1111111001111000001111111;
    rom[1091] = 25'b1111111001110101000000101;
    rom[1092] = 25'b1111111001110001111001000;
    rom[1093] = 25'b1111111001101110111000110;
    rom[1094] = 25'b1111111001101100000000001;
    rom[1095] = 25'b1111111001101001001111010;
    rom[1096] = 25'b1111111001100110100110001;
    rom[1097] = 25'b1111111001100100000101001;
    rom[1098] = 25'b1111111001100001101100001;
    rom[1099] = 25'b1111111001011111011011011;
    rom[1100] = 25'b1111111001011101010010111;
    rom[1101] = 25'b1111111001011011010010110;
    rom[1102] = 25'b1111111001011001011011001;
    rom[1103] = 25'b1111111001010111101100010;
    rom[1104] = 25'b1111111001010110000110000;
    rom[1105] = 25'b1111111001010100101000101;
    rom[1106] = 25'b1111111001010011010100001;
    rom[1107] = 25'b1111111001010010001000110;
    rom[1108] = 25'b1111111001010001000110011;
    rom[1109] = 25'b1111111001010000001101010;
    rom[1110] = 25'b1111111001001111011101010;
    rom[1111] = 25'b1111111001001110110110110;
    rom[1112] = 25'b1111111001001110011001110;
    rom[1113] = 25'b1111111001001110000110010;
    rom[1114] = 25'b1111111001001101111100010;
    rom[1115] = 25'b1111111001001101111100000;
    rom[1116] = 25'b1111111001001110000101011;
    rom[1117] = 25'b1111111001001110011000101;
    rom[1118] = 25'b1111111001001110110101110;
    rom[1119] = 25'b1111111001001111011100111;
    rom[1120] = 25'b1111111001010000001101111;
    rom[1121] = 25'b1111111001010001001001000;
    rom[1122] = 25'b1111111001010010001110001;
    rom[1123] = 25'b1111111001010011011101100;
    rom[1124] = 25'b1111111001010100110110111;
    rom[1125] = 25'b1111111001010110011010101;
    rom[1126] = 25'b1111111001011000001000101;
    rom[1127] = 25'b1111111001011010000000111;
    rom[1128] = 25'b1111111001011100000011100;
    rom[1129] = 25'b1111111001011110010000100;
    rom[1130] = 25'b1111111001100000100111111;
    rom[1131] = 25'b1111111001100011001001101;
    rom[1132] = 25'b1111111001100101110101110;
    rom[1133] = 25'b1111111001101000101100010;
    rom[1134] = 25'b1111111001101011101101011;
    rom[1135] = 25'b1111111001101110111000110;
    rom[1136] = 25'b1111111001110010001110101;
    rom[1137] = 25'b1111111001110101101111000;
    rom[1138] = 25'b1111111001111001011001111;
    rom[1139] = 25'b1111111001111101001111000;
    rom[1140] = 25'b1111111010000001001110101;
    rom[1141] = 25'b1111111010000101011000101;
    rom[1142] = 25'b1111111010001001101101001;
    rom[1143] = 25'b1111111010001110001011111;
    rom[1144] = 25'b1111111010010010110100111;
    rom[1145] = 25'b1111111010010111101000011;
    rom[1146] = 25'b1111111010011100100110000;
    rom[1147] = 25'b1111111010100001101101111;
    rom[1148] = 25'b1111111010100111000000000;
    rom[1149] = 25'b1111111010101100011100001;
    rom[1150] = 25'b1111111010110010000010011;
    rom[1151] = 25'b1111111010110111110010101;
    rom[1152] = 25'b1111111010111101101100111;
    rom[1153] = 25'b1111111011000011110001001;
    rom[1154] = 25'b1111111011001001111111001;
    rom[1155] = 25'b1111111011010000010110111;
    rom[1156] = 25'b1111111011010110111000010;
    rom[1157] = 25'b1111111011011101100011011;
    rom[1158] = 25'b1111111011100100010111111;
    rom[1159] = 25'b1111111011101011010110000;
    rom[1160] = 25'b1111111011110010011101011;
    rom[1161] = 25'b1111111011111001101101111;
    rom[1162] = 25'b1111111100000001000111110;
    rom[1163] = 25'b1111111100001000101010101;
    rom[1164] = 25'b1111111100010000010110010;
    rom[1165] = 25'b1111111100011000001011000;
    rom[1166] = 25'b1111111100100000001000010;
    rom[1167] = 25'b1111111100101000001110010;
    rom[1168] = 25'b1111111100110000011100101;
    rom[1169] = 25'b1111111100111000110011011;
    rom[1170] = 25'b1111111101000001010010011;
    rom[1171] = 25'b1111111101001001111001011;
    rom[1172] = 25'b1111111101010010101000011;
    rom[1173] = 25'b1111111101011011011111010;
    rom[1174] = 25'b1111111101100100011101110;
    rom[1175] = 25'b1111111101101101100011110;
    rom[1176] = 25'b1111111101110110110001001;
    rom[1177] = 25'b1111111110000000000101110;
    rom[1178] = 25'b1111111110001001100001011;
    rom[1179] = 25'b1111111110010011000011111;
    rom[1180] = 25'b1111111110011100101101001;
    rom[1181] = 25'b1111111110100110011100111;
    rom[1182] = 25'b1111111110110000010011000;
    rom[1183] = 25'b1111111110111010001111011;
    rom[1184] = 25'b1111111111000100010001110;
    rom[1185] = 25'b1111111111001110011001111;
    rom[1186] = 25'b1111111111011000100111110;
    rom[1187] = 25'b1111111111100010111011000;
    rom[1188] = 25'b1111111111101101010011101;
    rom[1189] = 25'b1111111111110111110001001;
    rom[1190] = 25'b0000000000000010010011101;
    rom[1191] = 25'b0000000000001100111010101;
    rom[1192] = 25'b0000000000010111100110010;
    rom[1193] = 25'b0000000000100010010110000;
    rom[1194] = 25'b0000000000101101001001111;
    rom[1195] = 25'b0000000000111000000001011;
    rom[1196] = 25'b0000000001000010111100101;
    rom[1197] = 25'b0000000001001101111011010;
    rom[1198] = 25'b0000000001011000111101000;
    rom[1199] = 25'b0000000001100100000001101;
    rom[1200] = 25'b0000000001101111001001000;
    rom[1201] = 25'b0000000001111010010010110;
    rom[1202] = 25'b0000000010000101011110111;
    rom[1203] = 25'b0000000010010000101100110;
    rom[1204] = 25'b0000000010011011111100101;
    rom[1205] = 25'b0000000010100111001101111;
    rom[1206] = 25'b0000000010110010100000011;
    rom[1207] = 25'b0000000010111101110100000;
    rom[1208] = 25'b0000000011001001001000010;
    rom[1209] = 25'b0000000011010100011101001;
    rom[1210] = 25'b0000000011011111110010010;
    rom[1211] = 25'b0000000011101011000111011;
    rom[1212] = 25'b0000000011110110011100010;
    rom[1213] = 25'b0000000100000001110000110;
    rom[1214] = 25'b0000000100001101000100011;
    rom[1215] = 25'b0000000100011000010111000;
    rom[1216] = 25'b0000000100100011101000011;
    rom[1217] = 25'b0000000100101110111000001;
    rom[1218] = 25'b0000000100111010000110010;
    rom[1219] = 25'b0000000101000101010010001;
    rom[1220] = 25'b0000000101010000011011110;
    rom[1221] = 25'b0000000101011011100010111;
    rom[1222] = 25'b0000000101100110100111000;
    rom[1223] = 25'b0000000101110001101000001;
    rom[1224] = 25'b0000000101111100100101110;
    rom[1225] = 25'b0000000110000111011111110;
    rom[1226] = 25'b0000000110010010010101110;
    rom[1227] = 25'b0000000110011101000111100;
    rom[1228] = 25'b0000000110100111110100111;
    rom[1229] = 25'b0000000110110010011101100;
    rom[1230] = 25'b0000000110111101000001001;
    rom[1231] = 25'b0000000111000111011111010;
    rom[1232] = 25'b0000000111010001111000000;
    rom[1233] = 25'b0000000111011100001010111;
    rom[1234] = 25'b0000000111100110010111101;
    rom[1235] = 25'b0000000111110000011110000;
    rom[1236] = 25'b0000000111111010011101101;
    rom[1237] = 25'b0000001000000100010110011;
    rom[1238] = 25'b0000001000001110000111111;
    rom[1239] = 25'b0000001000010111110010000;
    rom[1240] = 25'b0000001000100001010100011;
    rom[1241] = 25'b0000001000101010101110110;
    rom[1242] = 25'b0000001000110100000001000;
    rom[1243] = 25'b0000001000111101001010100;
    rom[1244] = 25'b0000001001000110001011011;
    rom[1245] = 25'b0000001001001111000011000;
    rom[1246] = 25'b0000001001010111110001100;
    rom[1247] = 25'b0000001001100000010110011;
    rom[1248] = 25'b0000001001101000110001011;
    rom[1249] = 25'b0000001001110001000010010;
    rom[1250] = 25'b0000001001111001001000110;
    rom[1251] = 25'b0000001010000001000100111;
    rom[1252] = 25'b0000001010001000110110000;
    rom[1253] = 25'b0000001010010000011100000;
    rom[1254] = 25'b0000001010010111110110110;
    rom[1255] = 25'b0000001010011111000101111;
    rom[1256] = 25'b0000001010100110001001010;
    rom[1257] = 25'b0000001010101101000000011;
    rom[1258] = 25'b0000001010110011101011011;
    rom[1259] = 25'b0000001010111010001001110;
    rom[1260] = 25'b0000001011000000011011011;
    rom[1261] = 25'b0000001011000110100000000;
    rom[1262] = 25'b0000001011001100010111100;
    rom[1263] = 25'b0000001011010010000001011;
    rom[1264] = 25'b0000001011010111011101110;
    rom[1265] = 25'b0000001011011100101100011;
    rom[1266] = 25'b0000001011100001101100110;
    rom[1267] = 25'b0000001011100110011110111;
    rom[1268] = 25'b0000001011101011000010011;
    rom[1269] = 25'b0000001011101111010111011;
    rom[1270] = 25'b0000001011110011011101100;
    rom[1271] = 25'b0000001011110111010100011;
    rom[1272] = 25'b0000001011111010111100001;
    rom[1273] = 25'b0000001011111110010100011;
    rom[1274] = 25'b0000001100000001011101000;
    rom[1275] = 25'b0000001100000100010101111;
    rom[1276] = 25'b0000001100000110111110101;
    rom[1277] = 25'b0000001100001001010111011;
    rom[1278] = 25'b0000001100001011011111110;
    rom[1279] = 25'b0000001100001101010111110;
    rom[1280] = 25'b0000001100001110111111000;
    rom[1281] = 25'b0000001100010000010101100;
    rom[1282] = 25'b0000001100010001011011001;
    rom[1283] = 25'b0000001100010010001111110;
    rom[1284] = 25'b0000001100010010110011001;
    rom[1285] = 25'b0000001100010011000101010;
    rom[1286] = 25'b0000001100010011000101111;
    rom[1287] = 25'b0000001100010010110101000;
    rom[1288] = 25'b0000001100010010010010100;
    rom[1289] = 25'b0000001100010001011110001;
    rom[1290] = 25'b0000001100010000011000000;
    rom[1291] = 25'b0000001100001110111111111;
    rom[1292] = 25'b0000001100001101010101101;
    rom[1293] = 25'b0000001100001011011001011;
    rom[1294] = 25'b0000001100001001001010110;
    rom[1295] = 25'b0000001100000110101001111;
    rom[1296] = 25'b0000001100000011110110110;
    rom[1297] = 25'b0000001100000000110001001;
    rom[1298] = 25'b0000001011111101011001000;
    rom[1299] = 25'b0000001011111001101110011;
    rom[1300] = 25'b0000001011110101110001011;
    rom[1301] = 25'b0000001011110001100001100;
    rom[1302] = 25'b0000001011101100111111001;
    rom[1303] = 25'b0000001011101000001010001;
    rom[1304] = 25'b0000001011100011000010100;
    rom[1305] = 25'b0000001011011101101000001;
    rom[1306] = 25'b0000001011010111111011001;
    rom[1307] = 25'b0000001011010001111011100;
    rom[1308] = 25'b0000001011001011101001000;
    rom[1309] = 25'b0000001011000101000100001;
    rom[1310] = 25'b0000001010111110001100011;
    rom[1311] = 25'b0000001010110111000010001;
    rom[1312] = 25'b0000001010101111100101011;
    rom[1313] = 25'b0000001010100111110110001;
    rom[1314] = 25'b0000001010011111110100010;
    rom[1315] = 25'b0000001010010111100000001;
    rom[1316] = 25'b0000001010001110111001100;
    rom[1317] = 25'b0000001010000110000000101;
    rom[1318] = 25'b0000001001111100110101101;
    rom[1319] = 25'b0000001001110011011000100;
    rom[1320] = 25'b0000001001101001101001011;
    rom[1321] = 25'b0000001001011111101000010;
    rom[1322] = 25'b0000001001010101010101011;
    rom[1323] = 25'b0000001001001010110000110;
    rom[1324] = 25'b0000001000111111111010011;
    rom[1325] = 25'b0000001000110100110010111;
    rom[1326] = 25'b0000001000101001011001110;
    rom[1327] = 25'b0000001000011101101111100;
    rom[1328] = 25'b0000001000010001110100010;
    rom[1329] = 25'b0000001000000101101000000;
    rom[1330] = 25'b0000000111111001001011001;
    rom[1331] = 25'b0000000111101100011101110;
    rom[1332] = 25'b0000000111011111011111110;
    rom[1333] = 25'b0000000111010010010001101;
    rom[1334] = 25'b0000000111000100110011100;
    rom[1335] = 25'b0000000110110111000101101;
    rom[1336] = 25'b0000000110101001001000000;
    rom[1337] = 25'b0000000110011010111011000;
    rom[1338] = 25'b0000000110001100011110110;
    rom[1339] = 25'b0000000101111101110011101;
    rom[1340] = 25'b0000000101101110111001101;
    rom[1341] = 25'b0000000101011111110001001;
    rom[1342] = 25'b0000000101010000011010010;
    rom[1343] = 25'b0000000101000000110101100;
    rom[1344] = 25'b0000000100110001000011000;
    rom[1345] = 25'b0000000100100001000010111;
    rom[1346] = 25'b0000000100010000110101100;
    rom[1347] = 25'b0000000100000000011011001;
    rom[1348] = 25'b0000000011101111110100010;
    rom[1349] = 25'b0000000011011111000000110;
    rom[1350] = 25'b0000000011001110000001010;
    rom[1351] = 25'b0000000010111100110101111;
    rom[1352] = 25'b0000000010101011011111000;
    rom[1353] = 25'b0000000010011001111101000;
    rom[1354] = 25'b0000000010001000010000000;
    rom[1355] = 25'b0000000001110110011000101;
    rom[1356] = 25'b0000000001100100010110111;
    rom[1357] = 25'b0000000001010010001011010;
    rom[1358] = 25'b0000000000111111110110000;
    rom[1359] = 25'b0000000000101101010111101;
    rom[1360] = 25'b0000000000011010110000011;
    rom[1361] = 25'b0000000000001000000000101;
    rom[1362] = 25'b1111111111110101001000111;
    rom[1363] = 25'b1111111111100010001001010;
    rom[1364] = 25'b1111111111001111000010010;
    rom[1365] = 25'b1111111110111011110100010;
    rom[1366] = 25'b1111111110101000011111100;
    rom[1367] = 25'b1111111110010101000100100;
    rom[1368] = 25'b1111111110000001100011110;
    rom[1369] = 25'b1111111101101101111101011;
    rom[1370] = 25'b1111111101011010010010001;
    rom[1371] = 25'b1111111101000110100010001;
    rom[1372] = 25'b1111111100110010101101111;
    rom[1373] = 25'b1111111100011110110101110;
    rom[1374] = 25'b1111111100001010111010011;
    rom[1375] = 25'b1111111011110110111011111;
    rom[1376] = 25'b1111111011100010111010110;
    rom[1377] = 25'b1111111011001110110111101;
    rom[1378] = 25'b1111111010111010110010110;
    rom[1379] = 25'b1111111010100110101100101;
    rom[1380] = 25'b1111111010010010100101101;
    rom[1381] = 25'b1111111001111110011110011;
    rom[1382] = 25'b1111111001101010010111000;
    rom[1383] = 25'b1111111001010110010000001;
    rom[1384] = 25'b1111111001000010001010011;
    rom[1385] = 25'b1111111000101110000101111;
    rom[1386] = 25'b1111111000011010000011011;
    rom[1387] = 25'b1111111000000110000011001;
    rom[1388] = 25'b1111110111110010000101101;
    rom[1389] = 25'b1111110111011110001011100;
    rom[1390] = 25'b1111110111001010010101000;
    rom[1391] = 25'b1111110110110110100010110;
    rom[1392] = 25'b1111110110100010110101000;
    rom[1393] = 25'b1111110110001111001100100;
    rom[1394] = 25'b1111110101111011101001101;
    rom[1395] = 25'b1111110101101000001100101;
    rom[1396] = 25'b1111110101010100110110011;
    rom[1397] = 25'b1111110101000001100111000;
    rom[1398] = 25'b1111110100101110011111001;
    rom[1399] = 25'b1111110100011011011111011;
    rom[1400] = 25'b1111110100001000100111111;
    rom[1401] = 25'b1111110011110101111001011;
    rom[1402] = 25'b1111110011100011010100001;
    rom[1403] = 25'b1111110011010000111000111;
    rom[1404] = 25'b1111110010111110100111111;
    rom[1405] = 25'b1111110010101100100001110;
    rom[1406] = 25'b1111110010011010100110111;
    rom[1407] = 25'b1111110010001000110111110;
    rom[1408] = 25'b1111110001110111010100111;
    rom[1409] = 25'b1111110001100101111110101;
    rom[1410] = 25'b1111110001010100110101101;
    rom[1411] = 25'b1111110001000011111010010;
    rom[1412] = 25'b1111110000110011001100111;
    rom[1413] = 25'b1111110000100010101110001;
    rom[1414] = 25'b1111110000010010011110100;
    rom[1415] = 25'b1111110000000010011110010;
    rom[1416] = 25'b1111101111110010101110000;
    rom[1417] = 25'b1111101111100011001110000;
    rom[1418] = 25'b1111101111010011111111000;
    rom[1419] = 25'b1111101111000101000001010;
    rom[1420] = 25'b1111101110110110010101010;
    rom[1421] = 25'b1111101110100111111011100;
    rom[1422] = 25'b1111101110011001110100010;
    rom[1423] = 25'b1111101110001100000000010;
    rom[1424] = 25'b1111101101111110011111101;
    rom[1425] = 25'b1111101101110001010010111;
    rom[1426] = 25'b1111101101100100011010100;
    rom[1427] = 25'b1111101101010111110111000;
    rom[1428] = 25'b1111101101001011101000100;
    rom[1429] = 25'b1111101100111111101111110;
    rom[1430] = 25'b1111101100110100001101000;
    rom[1431] = 25'b1111101100101001000000101;
    rom[1432] = 25'b1111101100011110001011000;
    rom[1433] = 25'b1111101100010011101100100;
    rom[1434] = 25'b1111101100001001100101101;
    rom[1435] = 25'b1111101011111111110110110;
    rom[1436] = 25'b1111101011110110100000001;
    rom[1437] = 25'b1111101011101101100010010;
    rom[1438] = 25'b1111101011100100111101011;
    rom[1439] = 25'b1111101011011100110010000;
    rom[1440] = 25'b1111101011010101000000010;
    rom[1441] = 25'b1111101011001101101000101;
    rom[1442] = 25'b1111101011000110101011100;
    rom[1443] = 25'b1111101011000000001001000;
    rom[1444] = 25'b1111101010111010000001110;
    rom[1445] = 25'b1111101010110100010101110;
    rom[1446] = 25'b1111101010101111000101100;
    rom[1447] = 25'b1111101010101010010001010;
    rom[1448] = 25'b1111101010100101111001010;
    rom[1449] = 25'b1111101010100001111101111;
    rom[1450] = 25'b1111101010011110011111010;
    rom[1451] = 25'b1111101010011011011101110;
    rom[1452] = 25'b1111101010011000111001101;
    rom[1453] = 25'b1111101010010110110011001;
    rom[1454] = 25'b1111101010010101001010101;
    rom[1455] = 25'b1111101010010100000000000;
    rom[1456] = 25'b1111101010010011010011111;
    rom[1457] = 25'b1111101010010011000110001;
    rom[1458] = 25'b1111101010010011010111001;
    rom[1459] = 25'b1111101010010100000111001;
    rom[1460] = 25'b1111101010010101010110010;
    rom[1461] = 25'b1111101010010111000100101;
    rom[1462] = 25'b1111101010011001010010011;
    rom[1463] = 25'b1111101010011011111111111;
    rom[1464] = 25'b1111101010011111001101000;
    rom[1465] = 25'b1111101010100010111010001;
    rom[1466] = 25'b1111101010100111000111010;
    rom[1467] = 25'b1111101010101011110100101;
    rom[1468] = 25'b1111101010110001000010001;
    rom[1469] = 25'b1111101010110110110000000;
    rom[1470] = 25'b1111101010111100111110010;
    rom[1471] = 25'b1111101011000011101101001;
    rom[1472] = 25'b1111101011001010111100100;
    rom[1473] = 25'b1111101011010010101100100;
    rom[1474] = 25'b1111101011011010111101010;
    rom[1475] = 25'b1111101011100011101110101;
    rom[1476] = 25'b1111101011101101000000110;
    rom[1477] = 25'b1111101011110110110011101;
    rom[1478] = 25'b1111101100000001000111010;
    rom[1479] = 25'b1111101100001011111011100;
    rom[1480] = 25'b1111101100010111010000101;
    rom[1481] = 25'b1111101100100011000110010;
    rom[1482] = 25'b1111101100101111011100100;
    rom[1483] = 25'b1111101100111100010011011;
    rom[1484] = 25'b1111101101001001101010110;
    rom[1485] = 25'b1111101101010111100010011;
    rom[1486] = 25'b1111101101100101111010100;
    rom[1487] = 25'b1111101101110100110010101;
    rom[1488] = 25'b1111101110000100001011000;
    rom[1489] = 25'b1111101110010100000011010;
    rom[1490] = 25'b1111101110100100011011011;
    rom[1491] = 25'b1111101110110101010011010;
    rom[1492] = 25'b1111101111000110101010011;
    rom[1493] = 25'b1111101111011000100001001;
    rom[1494] = 25'b1111101111101010110110111;
    rom[1495] = 25'b1111101111111101101011100;
    rom[1496] = 25'b1111110000010000111110111;
    rom[1497] = 25'b1111110000100100110000111;
    rom[1498] = 25'b1111110000111001000001000;
    rom[1499] = 25'b1111110001001101101111010;
    rom[1500] = 25'b1111110001100010111011001;
    rom[1501] = 25'b1111110001111000100100101;
    rom[1502] = 25'b1111110010001110101011010;
    rom[1503] = 25'b1111110010100101001110111;
    rom[1504] = 25'b1111110010111100001111000;
    rom[1505] = 25'b1111110011010011101011100;
    rom[1506] = 25'b1111110011101011100011111;
    rom[1507] = 25'b1111110100000011110111111;
    rom[1508] = 25'b1111110100011100100111010;
    rom[1509] = 25'b1111110100110101110001011;
    rom[1510] = 25'b1111110101001111010110001;
    rom[1511] = 25'b1111110101101001010100111;
    rom[1512] = 25'b1111110110000011101101100;
    rom[1513] = 25'b1111110110011110011111011;
    rom[1514] = 25'b1111110110111001101010001;
    rom[1515] = 25'b1111110111010101001101010;
    rom[1516] = 25'b1111110111110001001000100;
    rom[1517] = 25'b1111111000001101011011011;
    rom[1518] = 25'b1111111000101010000101001;
    rom[1519] = 25'b1111111001000111000101101;
    rom[1520] = 25'b1111111001100100011100010;
    rom[1521] = 25'b1111111010000010001000100;
    rom[1522] = 25'b1111111010100000001001111;
    rom[1523] = 25'b1111111010111110011111110;
    rom[1524] = 25'b1111111011011101001001110;
    rom[1525] = 25'b1111111011111100000111010;
    rom[1526] = 25'b1111111100011011010111101;
    rom[1527] = 25'b1111111100111010111010100;
    rom[1528] = 25'b1111111101011010101111010;
    rom[1529] = 25'b1111111101111010110101001;
    rom[1530] = 25'b1111111110011011001011110;
    rom[1531] = 25'b1111111110111011110010011;
    rom[1532] = 25'b1111111111011100101000100;
    rom[1533] = 25'b1111111111111101101101011;
    rom[1534] = 25'b0000000000011111000000011;
    rom[1535] = 25'b0000000001000000100001000;
    rom[1536] = 25'b0000000001100010001110100;
    rom[1537] = 25'b0000000010000100001000011;
    rom[1538] = 25'b0000000010100110001101110;
    rom[1539] = 25'b0000000011001000011110000;
    rom[1540] = 25'b0000000011101010111000101;
    rom[1541] = 25'b0000000100001101011100101;
    rom[1542] = 25'b0000000100110000001001101;
    rom[1543] = 25'b0000000101010010111110101;
    rom[1544] = 25'b0000000101110101111011001;
    rom[1545] = 25'b0000000110011000111110100;
    rom[1546] = 25'b0000000110111100000111101;
    rom[1547] = 25'b0000000111011111010110001;
    rom[1548] = 25'b0000001000000010101001001;
    rom[1549] = 25'b0000001000100101111111111;
    rom[1550] = 25'b0000001001001001011001101;
    rom[1551] = 25'b0000001001101100110101110;
    rom[1552] = 25'b0000001010010000010011010;
    rom[1553] = 25'b0000001010110011110001100;
    rom[1554] = 25'b0000001011010111001111110;
    rom[1555] = 25'b0000001011111010101101010;
    rom[1556] = 25'b0000001100011110001001000;
    rom[1557] = 25'b0000001101000001100010100;
    rom[1558] = 25'b0000001101100100111000110;
    rom[1559] = 25'b0000001110001000001011000;
    rom[1560] = 25'b0000001110101011011000100;
    rom[1561] = 25'b0000001111001110100000011;
    rom[1562] = 25'b0000001111110001100001111;
    rom[1563] = 25'b0000010000010100011100001;
    rom[1564] = 25'b0000010000110111001110011;
    rom[1565] = 25'b0000010001011001110111110;
    rom[1566] = 25'b0000010001111100010111101;
    rom[1567] = 25'b0000010010011110101100111;
    rom[1568] = 25'b0000010011000000110110111;
    rom[1569] = 25'b0000010011100010110100110;
    rom[1570] = 25'b0000010100000100100101101;
    rom[1571] = 25'b0000010100100110001000110;
    rom[1572] = 25'b0000010101000111011101010;
    rom[1573] = 25'b0000010101101000100010010;
    rom[1574] = 25'b0000010110001001010111001;
    rom[1575] = 25'b0000010110101001111010111;
    rom[1576] = 25'b0000010111001010001100101;
    rom[1577] = 25'b0000010111101010001011101;
    rom[1578] = 25'b0000011000001001110111000;
    rom[1579] = 25'b0000011000101001001110001;
    rom[1580] = 25'b0000011001001000001111111;
    rom[1581] = 25'b0000011001100110111011101;
    rom[1582] = 25'b0000011010000101010000100;
    rom[1583] = 25'b0000011010100011001101101;
    rom[1584] = 25'b0000011011000000110010011;
    rom[1585] = 25'b0000011011011101111101101;
    rom[1586] = 25'b0000011011111010101110110;
    rom[1587] = 25'b0000011100010111000101000;
    rom[1588] = 25'b0000011100110010111111100;
    rom[1589] = 25'b0000011101001110011101100;
    rom[1590] = 25'b0000011101101001011110001;
    rom[1591] = 25'b0000011110000100000000100;
    rom[1592] = 25'b0000011110011110000100000;
    rom[1593] = 25'b0000011110110111100111111;
    rom[1594] = 25'b0000011111010000101011010;
    rom[1595] = 25'b0000011111101001001101011;
    rom[1596] = 25'b0000100000000001001101011;
    rom[1597] = 25'b0000100000011000101010110;
    rom[1598] = 25'b0000100000101111100100100;
    rom[1599] = 25'b0000100001000101111010000;
    rom[1600] = 25'b0000100001011011101010101;
    rom[1601] = 25'b0000100001110000110101011;
    rom[1602] = 25'b0000100010000101011001110;
    rom[1603] = 25'b0000100010011001010111000;
    rom[1604] = 25'b0000100010101100101100010;
    rom[1605] = 25'b0000100010111111011001000;
    rom[1606] = 25'b0000100011010001011100011;
    rom[1607] = 25'b0000100011100010110110000;
    rom[1608] = 25'b0000100011110011100101000;
    rom[1609] = 25'b0000100100000011101000101;
    rom[1610] = 25'b0000100100010011000000011;
    rom[1611] = 25'b0000100100100001101011101;
    rom[1612] = 25'b0000100100101111101001101;
    rom[1613] = 25'b0000100100111100111001111;
    rom[1614] = 25'b0000100101001001011011110;
    rom[1615] = 25'b0000100101010101001110100;
    rom[1616] = 25'b0000100101100000010001110;
    rom[1617] = 25'b0000100101101010100100111;
    rom[1618] = 25'b0000100101110100000111010;
    rom[1619] = 25'b0000100101111100111000011;
    rom[1620] = 25'b0000100110000100110111101;
    rom[1621] = 25'b0000100110001100000100101;
    rom[1622] = 25'b0000100110010010011110110;
    rom[1623] = 25'b0000100110011000000101101;
    rom[1624] = 25'b0000100110011100111000101;
    rom[1625] = 25'b0000100110100000110111011;
    rom[1626] = 25'b0000100110100100000001100;
    rom[1627] = 25'b0000100110100110010110011;
    rom[1628] = 25'b0000100110100111110101101;
    rom[1629] = 25'b0000100110101000011110111;
    rom[1630] = 25'b0000100110101000010001111;
    rom[1631] = 25'b0000100110100111001101111;
    rom[1632] = 25'b0000100110100101010011000;
    rom[1633] = 25'b0000100110100010100000011;
    rom[1634] = 25'b0000100110011110110110001;
    rom[1635] = 25'b0000100110011010010011110;
    rom[1636] = 25'b0000100110010100111001000;
    rom[1637] = 25'b0000100110001110100101011;
    rom[1638] = 25'b0000100110000111011000111;
    rom[1639] = 25'b0000100101111111010011010;
    rom[1640] = 25'b0000100101110110010100000;
    rom[1641] = 25'b0000100101101100011011010;
    rom[1642] = 25'b0000100101100001101000100;
    rom[1643] = 25'b0000100101010101111011110;
    rom[1644] = 25'b0000100101001001010100111;
    rom[1645] = 25'b0000100100111011110011101;
    rom[1646] = 25'b0000100100101101010111111;
    rom[1647] = 25'b0000100100011110000001101;
    rom[1648] = 25'b0000100100001101110000110;
    rom[1649] = 25'b0000100011111100100101000;
    rom[1650] = 25'b0000100011101010011110101;
    rom[1651] = 25'b0000100011010111011101011;
    rom[1652] = 25'b0000100011000011100001011;
    rom[1653] = 25'b0000100010101110101010101;
    rom[1654] = 25'b0000100010011000111000111;
    rom[1655] = 25'b0000100010000010001100101;
    rom[1656] = 25'b0000100001101010100101101;
    rom[1657] = 25'b0000100001010010000100001;
    rom[1658] = 25'b0000100000111000101000001;
    rom[1659] = 25'b0000100000011110010001110;
    rom[1660] = 25'b0000100000000011000001001;
    rom[1661] = 25'b0000011111100110110110101;
    rom[1662] = 25'b0000011111001001110010010;
    rom[1663] = 25'b0000011110101011110100001;
    rom[1664] = 25'b0000011110001100111100101;
    rom[1665] = 25'b0000011101101101001100001;
    rom[1666] = 25'b0000011101001100100010100;
    rom[1667] = 25'b0000011100101011000000100;
    rom[1668] = 25'b0000011100001000100110001;
    rom[1669] = 25'b0000011011100101010011110;
    rom[1670] = 25'b0000011011000001001001111;
    rom[1671] = 25'b0000011010011100001000100;
    rom[1672] = 25'b0000011001110110010000100;
    rom[1673] = 25'b0000011001001111100010001;
    rom[1674] = 25'b0000011000100111111101101;
    rom[1675] = 25'b0000010111111111100011101;
    rom[1676] = 25'b0000010111010110010100100;
    rom[1677] = 25'b0000010110101100010000111;
    rom[1678] = 25'b0000010110000001011001001;
    rom[1679] = 25'b0000010101010101101101111;
    rom[1680] = 25'b0000010100101001001111101;
    rom[1681] = 25'b0000010011111011111111000;
    rom[1682] = 25'b0000010011001101111100101;
    rom[1683] = 25'b0000010010011111001001000;
    rom[1684] = 25'b0000010001101111100100111;
    rom[1685] = 25'b0000010000111111010000111;
    rom[1686] = 25'b0000010000001110001101101;
    rom[1687] = 25'b0000001111011100011100000;
    rom[1688] = 25'b0000001110101001111100100;
    rom[1689] = 25'b0000001101110110110000000;
    rom[1690] = 25'b0000001101000010110111001;
    rom[1691] = 25'b0000001100001110010010111;
    rom[1692] = 25'b0000001011011001000100000;
    rom[1693] = 25'b0000001010100011001011000;
    rom[1694] = 25'b0000001001101100101001010;
    rom[1695] = 25'b0000001000110101011111000;
    rom[1696] = 25'b0000000111111101101101101;
    rom[1697] = 25'b0000000111000101010101110;
    rom[1698] = 25'b0000000110001100011000100;
    rom[1699] = 25'b0000000101010010110110100;
    rom[1700] = 25'b0000000100011000110001001;
    rom[1701] = 25'b0000000011011110001000111;
    rom[1702] = 25'b0000000010100010111111000;
    rom[1703] = 25'b0000000001100111010100101;
    rom[1704] = 25'b0000000000101011001010100;
    rom[1705] = 25'b1111111111101110100001111;
    rom[1706] = 25'b1111111110110001011011101;
    rom[1707] = 25'b1111111101110011111001000;
    rom[1708] = 25'b1111111100110101111011000;
    rom[1709] = 25'b1111111011110111100010110;
    rom[1710] = 25'b1111111010111000110001010;
    rom[1711] = 25'b1111111001111001100111111;
    rom[1712] = 25'b1111111000111010000111110;
    rom[1713] = 25'b1111110111111010010001111;
    rom[1714] = 25'b1111110110111010000111101;
    rom[1715] = 25'b1111110101111001101010000;
    rom[1716] = 25'b1111110100111000111010100;
    rom[1717] = 25'b1111110011110111111010001;
    rom[1718] = 25'b1111110010110110101010011;
    rom[1719] = 25'b1111110001110101001100001;
    rom[1720] = 25'b1111110000110011100001000;
    rom[1721] = 25'b1111101111110001101010001;
    rom[1722] = 25'b1111101110101111101001000;
    rom[1723] = 25'b1111101101101101011110101;
    rom[1724] = 25'b1111101100101011001100100;
    rom[1725] = 25'b1111101011101000110100001;
    rom[1726] = 25'b1111101010100110010110101;
    rom[1727] = 25'b1111101001100011110101100;
    rom[1728] = 25'b1111101000100001010001111;
    rom[1729] = 25'b1111100111011110101101100;
    rom[1730] = 25'b1111100110011100001001110;
    rom[1731] = 25'b1111100101011001100111110;
    rom[1732] = 25'b1111100100010111001001001;
    rom[1733] = 25'b1111100011010100101111011;
    rom[1734] = 25'b1111100010010010011011101;
    rom[1735] = 25'b1111100001010000001111110;
    rom[1736] = 25'b1111100000001110001100111;
    rom[1737] = 25'b1111011111001100010100100;
    rom[1738] = 25'b1111011110001010101000010;
    rom[1739] = 25'b1111011101001001001001101;
    rom[1740] = 25'b1111011100000111111010000;
    rom[1741] = 25'b1111011011000110111011000;
    rom[1742] = 25'b1111011010000110001110000;
    rom[1743] = 25'b1111011001000101110100100;
    rom[1744] = 25'b1111011000000101110000001;
    rom[1745] = 25'b1111010111000110000010011;
    rom[1746] = 25'b1111010110000110101100101;
    rom[1747] = 25'b1111010101000111110000101;
    rom[1748] = 25'b1111010100001001001111110;
    rom[1749] = 25'b1111010011001011001011101;
    rom[1750] = 25'b1111010010001101100101110;
    rom[1751] = 25'b1111010001010000011111110;
    rom[1752] = 25'b1111010000010011111011000;
    rom[1753] = 25'b1111001111010111111001010;
    rom[1754] = 25'b1111001110011100011011111;
    rom[1755] = 25'b1111001101100001100100101;
    rom[1756] = 25'b1111001100100111010100111;
    rom[1757] = 25'b1111001011101101101110010;
    rom[1758] = 25'b1111001010110100110010010;
    rom[1759] = 25'b1111001001111100100010100;
    rom[1760] = 25'b1111001001000101000000100;
    rom[1761] = 25'b1111001000001110001101111;
    rom[1762] = 25'b1111000111011000001100000;
    rom[1763] = 25'b1111000110100010111100101;
    rom[1764] = 25'b1111000101101110100001010;
    rom[1765] = 25'b1111000100111010111011010;
    rom[1766] = 25'b1111000100001000001100011;
    rom[1767] = 25'b1111000011010110010110000;
    rom[1768] = 25'b1111000010100101011001110;
    rom[1769] = 25'b1111000001110101011001000;
    rom[1770] = 25'b1111000001000110010101100;
    rom[1771] = 25'b1111000000011000010000101;
    rom[1772] = 25'b1110111111101011001011111;
    rom[1773] = 25'b1110111110111111001000101;
    rom[1774] = 25'b1110111110010100001000101;
    rom[1775] = 25'b1110111101101010001101010;
    rom[1776] = 25'b1110111101000001010111110;
    rom[1777] = 25'b1110111100011001101010000;
    rom[1778] = 25'b1110111011110011000101001;
    rom[1779] = 25'b1110111011001101101010110;
    rom[1780] = 25'b1110111010101001011100010;
    rom[1781] = 25'b1110111010000110011011000;
    rom[1782] = 25'b1110111001100100101000100;
    rom[1783] = 25'b1110111001000100000110000;
    rom[1784] = 25'b1110111000100100110101001;
    rom[1785] = 25'b1110111000000110110111001;
    rom[1786] = 25'b1110110111101010001101011;
    rom[1787] = 25'b1110110111001110111001010;
    rom[1788] = 25'b1110110110110100111100000;
    rom[1789] = 25'b1110110110011100010111001;
    rom[1790] = 25'b1110110110000101001011101;
    rom[1791] = 25'b1110110101101111011011001;
    rom[1792] = 25'b1110110101011011000110110;
    rom[1793] = 25'b1110110101001000001111111;
    rom[1794] = 25'b1110110100110110110111101;
    rom[1795] = 25'b1110110100100110111111010;
    rom[1796] = 25'b1110110100011000100111111;
    rom[1797] = 25'b1110110100001011110011000;
    rom[1798] = 25'b1110110100000000100001101;
    rom[1799] = 25'b1110110011110110110100110;
    rom[1800] = 25'b1110110011101110101101110;
    rom[1801] = 25'b1110110011101000001101101;
    rom[1802] = 25'b1110110011100011010101101;
    rom[1803] = 25'b1110110011100000000110101;
    rom[1804] = 25'b1110110011011110100001110;
    rom[1805] = 25'b1110110011011110101000010;
    rom[1806] = 25'b1110110011100000011011000;
    rom[1807] = 25'b1110110011100011111010111;
    rom[1808] = 25'b1110110011101001001001000;
    rom[1809] = 25'b1110110011110000000110011;
    rom[1810] = 25'b1110110011111000110011110;
    rom[1811] = 25'b1110110100000011010010010;
    rom[1812] = 25'b1110110100001111100010101;
    rom[1813] = 25'b1110110100011101100101110;
    rom[1814] = 25'b1110110100101101011100101;
    rom[1815] = 25'b1110110100111111000111111;
    rom[1816] = 25'b1110110101010010101000011;
    rom[1817] = 25'b1110110101100111111110111;
    rom[1818] = 25'b1110110101111111001100000;
    rom[1819] = 25'b1110110110011000010000110;
    rom[1820] = 25'b1110110110110011001101101;
    rom[1821] = 25'b1110110111010000000011011;
    rom[1822] = 25'b1110110111101110110010100;
    rom[1823] = 25'b1110111000001111011011110;
    rom[1824] = 25'b1110111000110001111111101;
    rom[1825] = 25'b1110111001010110011110110;
    rom[1826] = 25'b1110111001111100111001101;
    rom[1827] = 25'b1110111010100101010000110;
    rom[1828] = 25'b1110111011001111100100110;
    rom[1829] = 25'b1110111011111011110101111;
    rom[1830] = 25'b1110111100101010000100100;
    rom[1831] = 25'b1110111101011010010001001;
    rom[1832] = 25'b1110111110001100011100001;
    rom[1833] = 25'b1110111111000000100110000;
    rom[1834] = 25'b1110111111110110101110101;
    rom[1835] = 25'b1111000000101110110110101;
    rom[1836] = 25'b1111000001101000111110001;
    rom[1837] = 25'b1111000010100101000101011;
    rom[1838] = 25'b1111000011100011001100100;
    rom[1839] = 25'b1111000100100011010011110;
    rom[1840] = 25'b1111000101100101011011001;
    rom[1841] = 25'b1111000110101001100010110;
    rom[1842] = 25'b1111000111101111101010110;
    rom[1843] = 25'b1111001000110111110011001;
    rom[1844] = 25'b1111001010000001111011111;
    rom[1845] = 25'b1111001011001110000100111;
    rom[1846] = 25'b1111001100011100001110010;
    rom[1847] = 25'b1111001101101100010111111;
    rom[1848] = 25'b1111001110111110100001100;
    rom[1849] = 25'b1111010000010010101010111;
    rom[1850] = 25'b1111010001101000110100000;
    rom[1851] = 25'b1111010011000000111100110;
    rom[1852] = 25'b1111010100011011000100101;
    rom[1853] = 25'b1111010101110111001011100;
    rom[1854] = 25'b1111010111010101010000111;
    rom[1855] = 25'b1111011000110101010100110;
    rom[1856] = 25'b1111011010010111010110011;
    rom[1857] = 25'b1111011011111011010101100;
    rom[1858] = 25'b1111011101100001010001101;
    rom[1859] = 25'b1111011111001001001010011;
    rom[1860] = 25'b1111100000110010111111001;
    rom[1861] = 25'b1111100010011110101111011;
    rom[1862] = 25'b1111100100001100011010101;
    rom[1863] = 25'b1111100101111100000000010;
    rom[1864] = 25'b1111100111101101011111011;
    rom[1865] = 25'b1111101001100000110111110;
    rom[1866] = 25'b1111101011010110001000011;
    rom[1867] = 25'b1111101101001101010000100;
    rom[1868] = 25'b1111101111000110001111100;
    rom[1869] = 25'b1111110001000001000100100;
    rom[1870] = 25'b1111110010111101101110110;
    rom[1871] = 25'b1111110100111100001101010;
    rom[1872] = 25'b1111110110111100011111010;
    rom[1873] = 25'b1111111000111110100011110;
    rom[1874] = 25'b1111111011000010011001110;
    rom[1875] = 25'b1111111101001000000000011;
    rom[1876] = 25'b1111111111001111010110101;
    rom[1877] = 25'b0000000001011000011011010;
    rom[1878] = 25'b0000000011100011001101011;
    rom[1879] = 25'b0000000101101111101011110;
    rom[1880] = 25'b0000000111111101110101011;
    rom[1881] = 25'b0000001010001101101001001;
    rom[1882] = 25'b0000001100011111000101101;
    rom[1883] = 25'b0000001110110010001001101;
    rom[1884] = 25'b0000010001000110110100000;
    rom[1885] = 25'b0000010011011101000011100;
    rom[1886] = 25'b0000010101110100110110101;
    rom[1887] = 25'b0000011000001110001100010;
    rom[1888] = 25'b0000011010101001000010110;
    rom[1889] = 25'b0000011101000101011001000;
    rom[1890] = 25'b0000011111100011001101011;
    rom[1891] = 25'b0000100010000010011110011;
    rom[1892] = 25'b0000100100100011001010101;
    rom[1893] = 25'b0000100111000101010000101;
    rom[1894] = 25'b0000101001101000101110110;
    rom[1895] = 25'b0000101100001101100011101;
    rom[1896] = 25'b0000101110110011101101100;
    rom[1897] = 25'b0000110001011011001010101;
    rom[1898] = 25'b0000110100000011111001101;
    rom[1899] = 25'b0000110110101101111000110;
    rom[1900] = 25'b0000111001011001000110001;
    rom[1901] = 25'b0000111100000101100000011;
    rom[1902] = 25'b0000111110110011000101011;
    rom[1903] = 25'b0001000001100001110011101;
    rom[1904] = 25'b0001000100010001101001010;
    rom[1905] = 25'b0001000111000010100100011;
    rom[1906] = 25'b0001001001110100100011010;
    rom[1907] = 25'b0001001100100111100100000;
    rom[1908] = 25'b0001001111011011100100110;
    rom[1909] = 25'b0001010010010000100011100;
    rom[1910] = 25'b0001010101000110011110011;
    rom[1911] = 25'b0001010111111101010011100;
    rom[1912] = 25'b0001011010110101000000111;
    rom[1913] = 25'b0001011101101101100100100;
    rom[1914] = 25'b0001100000100110111100010;
    rom[1915] = 25'b0001100011100001000110011;
    rom[1916] = 25'b0001100110011100000000101;
    rom[1917] = 25'b0001101001010111101001001;
    rom[1918] = 25'b0001101100010011111101100;
    rom[1919] = 25'b0001101111010000111011111;
    rom[1920] = 25'b0001110010001110100010001;
    rom[1921] = 25'b0001110101001100101101111;
    rom[1922] = 25'b0001111000001011011101011;
    rom[1923] = 25'b0001111011001010101110010;
    rom[1924] = 25'b0001111110001010011110011;
    rom[1925] = 25'b0010000001001010101011100;
    rom[1926] = 25'b0010000100001011010011011;
    rom[1927] = 25'b0010000111001100010011111;
    rom[1928] = 25'b0010001010001101101010111;
    rom[1929] = 25'b0010001101001111010110000;
    rom[1930] = 25'b0010010000010001010011000;
    rom[1931] = 25'b0010010011010011011111100;
    rom[1932] = 25'b0010010110010101111001100;
    rom[1933] = 25'b0010011001011000011110100;
    rom[1934] = 25'b0010011100011011001100011;
    rom[1935] = 25'b0010011111011110000000101;
    rom[1936] = 25'b0010100010100000111000111;
    rom[1937] = 25'b0010100101100011110011010;
    rom[1938] = 25'b0010101000100110101101000;
    rom[1939] = 25'b0010101011101001100011111;
    rom[1940] = 25'b0010101110101100010101101;
    rom[1941] = 25'b0010110001101110111111111;
    rom[1942] = 25'b0010110100110001100000010;
    rom[1943] = 25'b0010110111110011110100100;
    rom[1944] = 25'b0010111010110101111010000;
    rom[1945] = 25'b0010111101110111101110110;
    rom[1946] = 25'b0011000000111001010000001;
    rom[1947] = 25'b0011000011111010011011101;
    rom[1948] = 25'b0011000110111011001111010;
    rom[1949] = 25'b0011001001111011101000100;
    rom[1950] = 25'b0011001100111011100100111;
    rom[1951] = 25'b0011001111111011000010000;
    rom[1952] = 25'b0011010010111001111101101;
    rom[1953] = 25'b0011010101111000010101011;
    rom[1954] = 25'b0011011000110110000110111;
    rom[1955] = 25'b0011011011110011001111110;
    rom[1956] = 25'b0011011110101111101101100;
    rom[1957] = 25'b0011100001101011011110000;
    rom[1958] = 25'b0011100100100110011110101;
    rom[1959] = 25'b0011100111100000101101010;
    rom[1960] = 25'b0011101010011010000111011;
    rom[1961] = 25'b0011101101010010101010111;
    rom[1962] = 25'b0011110000001010010101001;
    rom[1963] = 25'b0011110011000001000100000;
    rom[1964] = 25'b0011110101110110110101001;
    rom[1965] = 25'b0011111000101011100110001;
    rom[1966] = 25'b0011111011011111010100110;
    rom[1967] = 25'b0011111110010001111110110;
    rom[1968] = 25'b0100000001000011100001111;
    rom[1969] = 25'b0100000011110011111011110;
    rom[1970] = 25'b0100000110100011001010001;
    rom[1971] = 25'b0100001001010001001010101;
    rom[1972] = 25'b0100001011111101111011010;
    rom[1973] = 25'b0100001110101001011001110;
    rom[1974] = 25'b0100010001010011100011110;
    rom[1975] = 25'b0100010011111100010111001;
    rom[1976] = 25'b0100010110100011110001101;
    rom[1977] = 25'b0100011001001001110001010;
    rom[1978] = 25'b0100011011101110010011110;
    rom[1979] = 25'b0100011110010001010110111;
    rom[1980] = 25'b0100100000110010111000110;
    rom[1981] = 25'b0100100011010010110111000;
    rom[1982] = 25'b0100100101110001001111110;
    rom[1983] = 25'b0100101000001110000000110;
    rom[1984] = 25'b0100101010101001001000001;
    rom[1985] = 25'b0100101101000010100011110;
    rom[1986] = 25'b0100101111011010010001100;
    rom[1987] = 25'b0100110001110000001111101;
    rom[1988] = 25'b0100110100000100011100000;
    rom[1989] = 25'b0100110110010110110100110;
    rom[1990] = 25'b0100111000100111010111111;
    rom[1991] = 25'b0100111010110110000011011;
    rom[1992] = 25'b0100111101000010110101101;
    rom[1993] = 25'b0100111111001101101100100;
    rom[1994] = 25'b0101000001010110100110011;
    rom[1995] = 25'b0101000011011101100001011;
    rom[1996] = 25'b0101000101100010011011101;
    rom[1997] = 25'b0101000111100101010011011;
    rom[1998] = 25'b0101001001100110000111000;
    rom[1999] = 25'b0101001011100100110100110;
    rom[2000] = 25'b0101001101100001011010110;
    rom[2001] = 25'b0101001111011011110111101;
    rom[2002] = 25'b0101010001010100001001101;
    rom[2003] = 25'b0101010011001010001111000;
    rom[2004] = 25'b0101010100111110000110011;
    rom[2005] = 25'b0101010110101111101110001;
    rom[2006] = 25'b0101011000011111000100111;
    rom[2007] = 25'b0101011010001100001000110;
    rom[2008] = 25'b0101011011110110111000110;
    rom[2009] = 25'b0101011101011111010011001;
    rom[2010] = 25'b0101011111000101010110110;
    rom[2011] = 25'b0101100000101001000001111;
    rom[2012] = 25'b0101100010001010010011011;
    rom[2013] = 25'b0101100011101001001010001;
    rom[2014] = 25'b0101100101000101100100100;
    rom[2015] = 25'b0101100110011111100001100;
    rom[2016] = 25'b0101100111110110111111111;
    rom[2017] = 25'b0101101001001011111110011;
    rom[2018] = 25'b0101101010011110011011111;
    rom[2019] = 25'b0101101011101110010111010;
    rom[2020] = 25'b0101101100111011101111100;
    rom[2021] = 25'b0101101110000110100011100;
    rom[2022] = 25'b0101101111001110110010010;
    rom[2023] = 25'b0101110000010100011010111;
    rom[2024] = 25'b0101110001010111011100011;
    rom[2025] = 25'b0101110010010111110101110;
    rom[2026] = 25'b0101110011010101100110010;
    rom[2027] = 25'b0101110100010000101101000;
    rom[2028] = 25'b0101110101001001001001001;
    rom[2029] = 25'b0101110101111110111010000;
    rom[2030] = 25'b0101110110110001111110110;
    rom[2031] = 25'b0101110111100010010110111;
    rom[2032] = 25'b0101111000010000000001100;
    rom[2033] = 25'b0101111000111010111110001;
    rom[2034] = 25'b0101111001100011001100001;
    rom[2035] = 25'b0101111010001000101011001;
    rom[2036] = 25'b0101111010101011011010011;
    rom[2037] = 25'b0101111011001011011001100;
    rom[2038] = 25'b0101111011101000101000001;
    rom[2039] = 25'b0101111100000011000101110;
    rom[2040] = 25'b0101111100011010110010000;
    rom[2041] = 25'b0101111100101111101100110;
    rom[2042] = 25'b0101111101000001110101100;
    rom[2043] = 25'b0101111101010001001100001;
    rom[2044] = 25'b0101111101011101110000011;
    rom[2045] = 25'b0101111101100111100010000;
    rom[2046] = 25'b0101111101101110100001000;
    rom[2047] = 25'b0101111101110010101101010;
    rom[2048] = 25'b0101111101110100000110110;
    rom[2049] = 25'b0101111101110010101101010;
    rom[2050] = 25'b0101111101101110100001000;
    rom[2051] = 25'b0101111101100111100010000;
    rom[2052] = 25'b0101111101011101110000011;
    rom[2053] = 25'b0101111101010001001100001;
    rom[2054] = 25'b0101111101000001110101100;
    rom[2055] = 25'b0101111100101111101100110;
    rom[2056] = 25'b0101111100011010110010000;
    rom[2057] = 25'b0101111100000011000101110;
    rom[2058] = 25'b0101111011101000101000001;
    rom[2059] = 25'b0101111011001011011001100;
    rom[2060] = 25'b0101111010101011011010011;
    rom[2061] = 25'b0101111010001000101011001;
    rom[2062] = 25'b0101111001100011001100001;
    rom[2063] = 25'b0101111000111010111110001;
    rom[2064] = 25'b0101111000010000000001100;
    rom[2065] = 25'b0101110111100010010110111;
    rom[2066] = 25'b0101110110110001111110110;
    rom[2067] = 25'b0101110101111110111010000;
    rom[2068] = 25'b0101110101001001001001001;
    rom[2069] = 25'b0101110100010000101101000;
    rom[2070] = 25'b0101110011010101100110010;
    rom[2071] = 25'b0101110010010111110101110;
    rom[2072] = 25'b0101110001010111011100011;
    rom[2073] = 25'b0101110000010100011010111;
    rom[2074] = 25'b0101101111001110110010010;
    rom[2075] = 25'b0101101110000110100011100;
    rom[2076] = 25'b0101101100111011101111100;
    rom[2077] = 25'b0101101011101110010111010;
    rom[2078] = 25'b0101101010011110011011111;
    rom[2079] = 25'b0101101001001011111110011;
    rom[2080] = 25'b0101100111110110111111111;
    rom[2081] = 25'b0101100110011111100001100;
    rom[2082] = 25'b0101100101000101100100100;
    rom[2083] = 25'b0101100011101001001010001;
    rom[2084] = 25'b0101100010001010010011011;
    rom[2085] = 25'b0101100000101001000001111;
    rom[2086] = 25'b0101011111000101010110110;
    rom[2087] = 25'b0101011101011111010011001;
    rom[2088] = 25'b0101011011110110111000110;
    rom[2089] = 25'b0101011010001100001000110;
    rom[2090] = 25'b0101011000011111000100111;
    rom[2091] = 25'b0101010110101111101110001;
    rom[2092] = 25'b0101010100111110000110011;
    rom[2093] = 25'b0101010011001010001111000;
    rom[2094] = 25'b0101010001010100001001101;
    rom[2095] = 25'b0101001111011011110111101;
    rom[2096] = 25'b0101001101100001011010110;
    rom[2097] = 25'b0101001011100100110100110;
    rom[2098] = 25'b0101001001100110000111000;
    rom[2099] = 25'b0101000111100101010011011;
    rom[2100] = 25'b0101000101100010011011101;
    rom[2101] = 25'b0101000011011101100001011;
    rom[2102] = 25'b0101000001010110100110011;
    rom[2103] = 25'b0100111111001101101100100;
    rom[2104] = 25'b0100111101000010110101101;
    rom[2105] = 25'b0100111010110110000011011;
    rom[2106] = 25'b0100111000100111010111111;
    rom[2107] = 25'b0100110110010110110100110;
    rom[2108] = 25'b0100110100000100011100000;
    rom[2109] = 25'b0100110001110000001111101;
    rom[2110] = 25'b0100101111011010010001100;
    rom[2111] = 25'b0100101101000010100011110;
    rom[2112] = 25'b0100101010101001001000001;
    rom[2113] = 25'b0100101000001110000000110;
    rom[2114] = 25'b0100100101110001001111110;
    rom[2115] = 25'b0100100011010010110111000;
    rom[2116] = 25'b0100100000110010111000110;
    rom[2117] = 25'b0100011110010001010110111;
    rom[2118] = 25'b0100011011101110010011110;
    rom[2119] = 25'b0100011001001001110001010;
    rom[2120] = 25'b0100010110100011110001101;
    rom[2121] = 25'b0100010011111100010111001;
    rom[2122] = 25'b0100010001010011100011110;
    rom[2123] = 25'b0100001110101001011001110;
    rom[2124] = 25'b0100001011111101111011010;
    rom[2125] = 25'b0100001001010001001010101;
    rom[2126] = 25'b0100000110100011001010001;
    rom[2127] = 25'b0100000011110011111011110;
    rom[2128] = 25'b0100000001000011100001111;
    rom[2129] = 25'b0011111110010001111110110;
    rom[2130] = 25'b0011111011011111010100110;
    rom[2131] = 25'b0011111000101011100110001;
    rom[2132] = 25'b0011110101110110110101001;
    rom[2133] = 25'b0011110011000001000100000;
    rom[2134] = 25'b0011110000001010010101001;
    rom[2135] = 25'b0011101101010010101010111;
    rom[2136] = 25'b0011101010011010000111011;
    rom[2137] = 25'b0011100111100000101101010;
    rom[2138] = 25'b0011100100100110011110101;
    rom[2139] = 25'b0011100001101011011110000;
    rom[2140] = 25'b0011011110101111101101100;
    rom[2141] = 25'b0011011011110011001111110;
    rom[2142] = 25'b0011011000110110000110111;
    rom[2143] = 25'b0011010101111000010101011;
    rom[2144] = 25'b0011010010111001111101101;
    rom[2145] = 25'b0011001111111011000010000;
    rom[2146] = 25'b0011001100111011100100111;
    rom[2147] = 25'b0011001001111011101000100;
    rom[2148] = 25'b0011000110111011001111010;
    rom[2149] = 25'b0011000011111010011011101;
    rom[2150] = 25'b0011000000111001010000001;
    rom[2151] = 25'b0010111101110111101110110;
    rom[2152] = 25'b0010111010110101111010000;
    rom[2153] = 25'b0010110111110011110100100;
    rom[2154] = 25'b0010110100110001100000010;
    rom[2155] = 25'b0010110001101110111111111;
    rom[2156] = 25'b0010101110101100010101101;
    rom[2157] = 25'b0010101011101001100011111;
    rom[2158] = 25'b0010101000100110101101000;
    rom[2159] = 25'b0010100101100011110011010;
    rom[2160] = 25'b0010100010100000111000111;
    rom[2161] = 25'b0010011111011110000000101;
    rom[2162] = 25'b0010011100011011001100011;
    rom[2163] = 25'b0010011001011000011110100;
    rom[2164] = 25'b0010010110010101111001100;
    rom[2165] = 25'b0010010011010011011111100;
    rom[2166] = 25'b0010010000010001010011000;
    rom[2167] = 25'b0010001101001111010110000;
    rom[2168] = 25'b0010001010001101101010111;
    rom[2169] = 25'b0010000111001100010011111;
    rom[2170] = 25'b0010000100001011010011011;
    rom[2171] = 25'b0010000001001010101011100;
    rom[2172] = 25'b0001111110001010011110011;
    rom[2173] = 25'b0001111011001010101110010;
    rom[2174] = 25'b0001111000001011011101011;
    rom[2175] = 25'b0001110101001100101101111;
    rom[2176] = 25'b0001110010001110100010001;
    rom[2177] = 25'b0001101111010000111011111;
    rom[2178] = 25'b0001101100010011111101100;
    rom[2179] = 25'b0001101001010111101001001;
    rom[2180] = 25'b0001100110011100000000101;
    rom[2181] = 25'b0001100011100001000110011;
    rom[2182] = 25'b0001100000100110111100010;
    rom[2183] = 25'b0001011101101101100100100;
    rom[2184] = 25'b0001011010110101000000111;
    rom[2185] = 25'b0001010111111101010011100;
    rom[2186] = 25'b0001010101000110011110011;
    rom[2187] = 25'b0001010010010000100011100;
    rom[2188] = 25'b0001001111011011100100110;
    rom[2189] = 25'b0001001100100111100100000;
    rom[2190] = 25'b0001001001110100100011010;
    rom[2191] = 25'b0001000111000010100100011;
    rom[2192] = 25'b0001000100010001101001010;
    rom[2193] = 25'b0001000001100001110011101;
    rom[2194] = 25'b0000111110110011000101011;
    rom[2195] = 25'b0000111100000101100000011;
    rom[2196] = 25'b0000111001011001000110001;
    rom[2197] = 25'b0000110110101101111000110;
    rom[2198] = 25'b0000110100000011111001101;
    rom[2199] = 25'b0000110001011011001010101;
    rom[2200] = 25'b0000101110110011101101100;
    rom[2201] = 25'b0000101100001101100011101;
    rom[2202] = 25'b0000101001101000101110110;
    rom[2203] = 25'b0000100111000101010000101;
    rom[2204] = 25'b0000100100100011001010101;
    rom[2205] = 25'b0000100010000010011110011;
    rom[2206] = 25'b0000011111100011001101011;
    rom[2207] = 25'b0000011101000101011001000;
    rom[2208] = 25'b0000011010101001000010110;
    rom[2209] = 25'b0000011000001110001100010;
    rom[2210] = 25'b0000010101110100110110101;
    rom[2211] = 25'b0000010011011101000011100;
    rom[2212] = 25'b0000010001000110110100000;
    rom[2213] = 25'b0000001110110010001001101;
    rom[2214] = 25'b0000001100011111000101101;
    rom[2215] = 25'b0000001010001101101001001;
    rom[2216] = 25'b0000000111111101110101011;
    rom[2217] = 25'b0000000101101111101011110;
    rom[2218] = 25'b0000000011100011001101011;
    rom[2219] = 25'b0000000001011000011011010;
    rom[2220] = 25'b1111111111001111010110101;
    rom[2221] = 25'b1111111101001000000000011;
    rom[2222] = 25'b1111111011000010011001110;
    rom[2223] = 25'b1111111000111110100011110;
    rom[2224] = 25'b1111110110111100011111010;
    rom[2225] = 25'b1111110100111100001101010;
    rom[2226] = 25'b1111110010111101101110110;
    rom[2227] = 25'b1111110001000001000100100;
    rom[2228] = 25'b1111101111000110001111100;
    rom[2229] = 25'b1111101101001101010000100;
    rom[2230] = 25'b1111101011010110001000011;
    rom[2231] = 25'b1111101001100000110111110;
    rom[2232] = 25'b1111100111101101011111011;
    rom[2233] = 25'b1111100101111100000000010;
    rom[2234] = 25'b1111100100001100011010101;
    rom[2235] = 25'b1111100010011110101111011;
    rom[2236] = 25'b1111100000110010111111001;
    rom[2237] = 25'b1111011111001001001010011;
    rom[2238] = 25'b1111011101100001010001101;
    rom[2239] = 25'b1111011011111011010101100;
    rom[2240] = 25'b1111011010010111010110011;
    rom[2241] = 25'b1111011000110101010100110;
    rom[2242] = 25'b1111010111010101010000111;
    rom[2243] = 25'b1111010101110111001011100;
    rom[2244] = 25'b1111010100011011000100101;
    rom[2245] = 25'b1111010011000000111100110;
    rom[2246] = 25'b1111010001101000110100000;
    rom[2247] = 25'b1111010000010010101010111;
    rom[2248] = 25'b1111001110111110100001100;
    rom[2249] = 25'b1111001101101100010111111;
    rom[2250] = 25'b1111001100011100001110010;
    rom[2251] = 25'b1111001011001110000100111;
    rom[2252] = 25'b1111001010000001111011111;
    rom[2253] = 25'b1111001000110111110011001;
    rom[2254] = 25'b1111000111101111101010110;
    rom[2255] = 25'b1111000110101001100010110;
    rom[2256] = 25'b1111000101100101011011001;
    rom[2257] = 25'b1111000100100011010011110;
    rom[2258] = 25'b1111000011100011001100100;
    rom[2259] = 25'b1111000010100101000101011;
    rom[2260] = 25'b1111000001101000111110001;
    rom[2261] = 25'b1111000000101110110110101;
    rom[2262] = 25'b1110111111110110101110101;
    rom[2263] = 25'b1110111111000000100110000;
    rom[2264] = 25'b1110111110001100011100001;
    rom[2265] = 25'b1110111101011010010001001;
    rom[2266] = 25'b1110111100101010000100100;
    rom[2267] = 25'b1110111011111011110101111;
    rom[2268] = 25'b1110111011001111100100110;
    rom[2269] = 25'b1110111010100101010000110;
    rom[2270] = 25'b1110111001111100111001101;
    rom[2271] = 25'b1110111001010110011110110;
    rom[2272] = 25'b1110111000110001111111101;
    rom[2273] = 25'b1110111000001111011011110;
    rom[2274] = 25'b1110110111101110110010100;
    rom[2275] = 25'b1110110111010000000011011;
    rom[2276] = 25'b1110110110110011001101101;
    rom[2277] = 25'b1110110110011000010000110;
    rom[2278] = 25'b1110110101111111001100000;
    rom[2279] = 25'b1110110101100111111110111;
    rom[2280] = 25'b1110110101010010101000011;
    rom[2281] = 25'b1110110100111111000111111;
    rom[2282] = 25'b1110110100101101011100101;
    rom[2283] = 25'b1110110100011101100101110;
    rom[2284] = 25'b1110110100001111100010101;
    rom[2285] = 25'b1110110100000011010010010;
    rom[2286] = 25'b1110110011111000110011110;
    rom[2287] = 25'b1110110011110000000110011;
    rom[2288] = 25'b1110110011101001001001000;
    rom[2289] = 25'b1110110011100011111010111;
    rom[2290] = 25'b1110110011100000011011000;
    rom[2291] = 25'b1110110011011110101000010;
    rom[2292] = 25'b1110110011011110100001110;
    rom[2293] = 25'b1110110011100000000110101;
    rom[2294] = 25'b1110110011100011010101101;
    rom[2295] = 25'b1110110011101000001101101;
    rom[2296] = 25'b1110110011101110101101110;
    rom[2297] = 25'b1110110011110110110100110;
    rom[2298] = 25'b1110110100000000100001101;
    rom[2299] = 25'b1110110100001011110011000;
    rom[2300] = 25'b1110110100011000100111111;
    rom[2301] = 25'b1110110100100110111111010;
    rom[2302] = 25'b1110110100110110110111101;
    rom[2303] = 25'b1110110101001000001111111;
    rom[2304] = 25'b1110110101011011000110110;
    rom[2305] = 25'b1110110101101111011011001;
    rom[2306] = 25'b1110110110000101001011101;
    rom[2307] = 25'b1110110110011100010111001;
    rom[2308] = 25'b1110110110110100111100000;
    rom[2309] = 25'b1110110111001110111001010;
    rom[2310] = 25'b1110110111101010001101011;
    rom[2311] = 25'b1110111000000110110111001;
    rom[2312] = 25'b1110111000100100110101001;
    rom[2313] = 25'b1110111001000100000110000;
    rom[2314] = 25'b1110111001100100101000100;
    rom[2315] = 25'b1110111010000110011011000;
    rom[2316] = 25'b1110111010101001011100010;
    rom[2317] = 25'b1110111011001101101010110;
    rom[2318] = 25'b1110111011110011000101001;
    rom[2319] = 25'b1110111100011001101010000;
    rom[2320] = 25'b1110111101000001010111110;
    rom[2321] = 25'b1110111101101010001101010;
    rom[2322] = 25'b1110111110010100001000101;
    rom[2323] = 25'b1110111110111111001000101;
    rom[2324] = 25'b1110111111101011001011111;
    rom[2325] = 25'b1111000000011000010000101;
    rom[2326] = 25'b1111000001000110010101100;
    rom[2327] = 25'b1111000001110101011001000;
    rom[2328] = 25'b1111000010100101011001110;
    rom[2329] = 25'b1111000011010110010110000;
    rom[2330] = 25'b1111000100001000001100011;
    rom[2331] = 25'b1111000100111010111011010;
    rom[2332] = 25'b1111000101101110100001010;
    rom[2333] = 25'b1111000110100010111100101;
    rom[2334] = 25'b1111000111011000001100000;
    rom[2335] = 25'b1111001000001110001101111;
    rom[2336] = 25'b1111001001000101000000100;
    rom[2337] = 25'b1111001001111100100010100;
    rom[2338] = 25'b1111001010110100110010010;
    rom[2339] = 25'b1111001011101101101110010;
    rom[2340] = 25'b1111001100100111010100111;
    rom[2341] = 25'b1111001101100001100100101;
    rom[2342] = 25'b1111001110011100011011111;
    rom[2343] = 25'b1111001111010111111001010;
    rom[2344] = 25'b1111010000010011111011000;
    rom[2345] = 25'b1111010001010000011111110;
    rom[2346] = 25'b1111010010001101100101110;
    rom[2347] = 25'b1111010011001011001011101;
    rom[2348] = 25'b1111010100001001001111110;
    rom[2349] = 25'b1111010101000111110000101;
    rom[2350] = 25'b1111010110000110101100101;
    rom[2351] = 25'b1111010111000110000010011;
    rom[2352] = 25'b1111011000000101110000001;
    rom[2353] = 25'b1111011001000101110100100;
    rom[2354] = 25'b1111011010000110001110000;
    rom[2355] = 25'b1111011011000110111011000;
    rom[2356] = 25'b1111011100000111111010000;
    rom[2357] = 25'b1111011101001001001001101;
    rom[2358] = 25'b1111011110001010101000010;
    rom[2359] = 25'b1111011111001100010100100;
    rom[2360] = 25'b1111100000001110001100111;
    rom[2361] = 25'b1111100001010000001111110;
    rom[2362] = 25'b1111100010010010011011101;
    rom[2363] = 25'b1111100011010100101111011;
    rom[2364] = 25'b1111100100010111001001001;
    rom[2365] = 25'b1111100101011001100111110;
    rom[2366] = 25'b1111100110011100001001110;
    rom[2367] = 25'b1111100111011110101101100;
    rom[2368] = 25'b1111101000100001010001111;
    rom[2369] = 25'b1111101001100011110101100;
    rom[2370] = 25'b1111101010100110010110101;
    rom[2371] = 25'b1111101011101000110100001;
    rom[2372] = 25'b1111101100101011001100100;
    rom[2373] = 25'b1111101101101101011110101;
    rom[2374] = 25'b1111101110101111101001000;
    rom[2375] = 25'b1111101111110001101010001;
    rom[2376] = 25'b1111110000110011100001000;
    rom[2377] = 25'b1111110001110101001100001;
    rom[2378] = 25'b1111110010110110101010011;
    rom[2379] = 25'b1111110011110111111010001;
    rom[2380] = 25'b1111110100111000111010100;
    rom[2381] = 25'b1111110101111001101010000;
    rom[2382] = 25'b1111110110111010000111101;
    rom[2383] = 25'b1111110111111010010001111;
    rom[2384] = 25'b1111111000111010000111110;
    rom[2385] = 25'b1111111001111001100111111;
    rom[2386] = 25'b1111111010111000110001010;
    rom[2387] = 25'b1111111011110111100010110;
    rom[2388] = 25'b1111111100110101111011000;
    rom[2389] = 25'b1111111101110011111001000;
    rom[2390] = 25'b1111111110110001011011101;
    rom[2391] = 25'b1111111111101110100001111;
    rom[2392] = 25'b0000000000101011001010100;
    rom[2393] = 25'b0000000001100111010100101;
    rom[2394] = 25'b0000000010100010111111000;
    rom[2395] = 25'b0000000011011110001000111;
    rom[2396] = 25'b0000000100011000110001001;
    rom[2397] = 25'b0000000101010010110110100;
    rom[2398] = 25'b0000000110001100011000100;
    rom[2399] = 25'b0000000111000101010101110;
    rom[2400] = 25'b0000000111111101101101101;
    rom[2401] = 25'b0000001000110101011111000;
    rom[2402] = 25'b0000001001101100101001010;
    rom[2403] = 25'b0000001010100011001011000;
    rom[2404] = 25'b0000001011011001000100000;
    rom[2405] = 25'b0000001100001110010010111;
    rom[2406] = 25'b0000001101000010110111001;
    rom[2407] = 25'b0000001101110110110000000;
    rom[2408] = 25'b0000001110101001111100100;
    rom[2409] = 25'b0000001111011100011100000;
    rom[2410] = 25'b0000010000001110001101101;
    rom[2411] = 25'b0000010000111111010000111;
    rom[2412] = 25'b0000010001101111100100111;
    rom[2413] = 25'b0000010010011111001001000;
    rom[2414] = 25'b0000010011001101111100101;
    rom[2415] = 25'b0000010011111011111111000;
    rom[2416] = 25'b0000010100101001001111101;
    rom[2417] = 25'b0000010101010101101101111;
    rom[2418] = 25'b0000010110000001011001001;
    rom[2419] = 25'b0000010110101100010000111;
    rom[2420] = 25'b0000010111010110010100100;
    rom[2421] = 25'b0000010111111111100011101;
    rom[2422] = 25'b0000011000100111111101101;
    rom[2423] = 25'b0000011001001111100010001;
    rom[2424] = 25'b0000011001110110010000100;
    rom[2425] = 25'b0000011010011100001000100;
    rom[2426] = 25'b0000011011000001001001111;
    rom[2427] = 25'b0000011011100101010011110;
    rom[2428] = 25'b0000011100001000100110001;
    rom[2429] = 25'b0000011100101011000000100;
    rom[2430] = 25'b0000011101001100100010100;
    rom[2431] = 25'b0000011101101101001100001;
    rom[2432] = 25'b0000011110001100111100101;
    rom[2433] = 25'b0000011110101011110100001;
    rom[2434] = 25'b0000011111001001110010010;
    rom[2435] = 25'b0000011111100110110110101;
    rom[2436] = 25'b0000100000000011000001001;
    rom[2437] = 25'b0000100000011110010001110;
    rom[2438] = 25'b0000100000111000101000001;
    rom[2439] = 25'b0000100001010010000100001;
    rom[2440] = 25'b0000100001101010100101101;
    rom[2441] = 25'b0000100010000010001100101;
    rom[2442] = 25'b0000100010011000111000111;
    rom[2443] = 25'b0000100010101110101010101;
    rom[2444] = 25'b0000100011000011100001011;
    rom[2445] = 25'b0000100011010111011101011;
    rom[2446] = 25'b0000100011101010011110101;
    rom[2447] = 25'b0000100011111100100101000;
    rom[2448] = 25'b0000100100001101110000110;
    rom[2449] = 25'b0000100100011110000001101;
    rom[2450] = 25'b0000100100101101010111111;
    rom[2451] = 25'b0000100100111011110011101;
    rom[2452] = 25'b0000100101001001010100111;
    rom[2453] = 25'b0000100101010101111011110;
    rom[2454] = 25'b0000100101100001101000100;
    rom[2455] = 25'b0000100101101100011011010;
    rom[2456] = 25'b0000100101110110010100000;
    rom[2457] = 25'b0000100101111111010011010;
    rom[2458] = 25'b0000100110000111011000111;
    rom[2459] = 25'b0000100110001110100101011;
    rom[2460] = 25'b0000100110010100111001000;
    rom[2461] = 25'b0000100110011010010011110;
    rom[2462] = 25'b0000100110011110110110001;
    rom[2463] = 25'b0000100110100010100000011;
    rom[2464] = 25'b0000100110100101010011000;
    rom[2465] = 25'b0000100110100111001101111;
    rom[2466] = 25'b0000100110101000010001111;
    rom[2467] = 25'b0000100110101000011110111;
    rom[2468] = 25'b0000100110100111110101101;
    rom[2469] = 25'b0000100110100110010110011;
    rom[2470] = 25'b0000100110100100000001100;
    rom[2471] = 25'b0000100110100000110111011;
    rom[2472] = 25'b0000100110011100111000101;
    rom[2473] = 25'b0000100110011000000101101;
    rom[2474] = 25'b0000100110010010011110110;
    rom[2475] = 25'b0000100110001100000100101;
    rom[2476] = 25'b0000100110000100110111101;
    rom[2477] = 25'b0000100101111100111000011;
    rom[2478] = 25'b0000100101110100000111010;
    rom[2479] = 25'b0000100101101010100100111;
    rom[2480] = 25'b0000100101100000010001110;
    rom[2481] = 25'b0000100101010101001110100;
    rom[2482] = 25'b0000100101001001011011110;
    rom[2483] = 25'b0000100100111100111001111;
    rom[2484] = 25'b0000100100101111101001101;
    rom[2485] = 25'b0000100100100001101011101;
    rom[2486] = 25'b0000100100010011000000011;
    rom[2487] = 25'b0000100100000011101000101;
    rom[2488] = 25'b0000100011110011100101000;
    rom[2489] = 25'b0000100011100010110110000;
    rom[2490] = 25'b0000100011010001011100011;
    rom[2491] = 25'b0000100010111111011001000;
    rom[2492] = 25'b0000100010101100101100010;
    rom[2493] = 25'b0000100010011001010111000;
    rom[2494] = 25'b0000100010000101011001110;
    rom[2495] = 25'b0000100001110000110101011;
    rom[2496] = 25'b0000100001011011101010101;
    rom[2497] = 25'b0000100001000101111010000;
    rom[2498] = 25'b0000100000101111100100100;
    rom[2499] = 25'b0000100000011000101010110;
    rom[2500] = 25'b0000100000000001001101011;
    rom[2501] = 25'b0000011111101001001101011;
    rom[2502] = 25'b0000011111010000101011010;
    rom[2503] = 25'b0000011110110111100111111;
    rom[2504] = 25'b0000011110011110000100000;
    rom[2505] = 25'b0000011110000100000000100;
    rom[2506] = 25'b0000011101101001011110001;
    rom[2507] = 25'b0000011101001110011101100;
    rom[2508] = 25'b0000011100110010111111100;
    rom[2509] = 25'b0000011100010111000101000;
    rom[2510] = 25'b0000011011111010101110110;
    rom[2511] = 25'b0000011011011101111101101;
    rom[2512] = 25'b0000011011000000110010011;
    rom[2513] = 25'b0000011010100011001101101;
    rom[2514] = 25'b0000011010000101010000100;
    rom[2515] = 25'b0000011001100110111011101;
    rom[2516] = 25'b0000011001001000001111111;
    rom[2517] = 25'b0000011000101001001110001;
    rom[2518] = 25'b0000011000001001110111000;
    rom[2519] = 25'b0000010111101010001011101;
    rom[2520] = 25'b0000010111001010001100101;
    rom[2521] = 25'b0000010110101001111010111;
    rom[2522] = 25'b0000010110001001010111001;
    rom[2523] = 25'b0000010101101000100010010;
    rom[2524] = 25'b0000010101000111011101010;
    rom[2525] = 25'b0000010100100110001000110;
    rom[2526] = 25'b0000010100000100100101101;
    rom[2527] = 25'b0000010011100010110100110;
    rom[2528] = 25'b0000010011000000110110111;
    rom[2529] = 25'b0000010010011110101100111;
    rom[2530] = 25'b0000010001111100010111101;
    rom[2531] = 25'b0000010001011001110111110;
    rom[2532] = 25'b0000010000110111001110011;
    rom[2533] = 25'b0000010000010100011100001;
    rom[2534] = 25'b0000001111110001100001111;
    rom[2535] = 25'b0000001111001110100000011;
    rom[2536] = 25'b0000001110101011011000100;
    rom[2537] = 25'b0000001110001000001011000;
    rom[2538] = 25'b0000001101100100111000110;
    rom[2539] = 25'b0000001101000001100010100;
    rom[2540] = 25'b0000001100011110001001000;
    rom[2541] = 25'b0000001011111010101101010;
    rom[2542] = 25'b0000001011010111001111110;
    rom[2543] = 25'b0000001010110011110001100;
    rom[2544] = 25'b0000001010010000010011010;
    rom[2545] = 25'b0000001001101100110101110;
    rom[2546] = 25'b0000001001001001011001101;
    rom[2547] = 25'b0000001000100101111111111;
    rom[2548] = 25'b0000001000000010101001001;
    rom[2549] = 25'b0000000111011111010110001;
    rom[2550] = 25'b0000000110111100000111101;
    rom[2551] = 25'b0000000110011000111110100;
    rom[2552] = 25'b0000000101110101111011001;
    rom[2553] = 25'b0000000101010010111110101;
    rom[2554] = 25'b0000000100110000001001101;
    rom[2555] = 25'b0000000100001101011100101;
    rom[2556] = 25'b0000000011101010111000101;
    rom[2557] = 25'b0000000011001000011110000;
    rom[2558] = 25'b0000000010100110001101110;
    rom[2559] = 25'b0000000010000100001000011;
    rom[2560] = 25'b0000000001100010001110100;
    rom[2561] = 25'b0000000001000000100001000;
    rom[2562] = 25'b0000000000011111000000011;
    rom[2563] = 25'b1111111111111101101101011;
    rom[2564] = 25'b1111111111011100101000100;
    rom[2565] = 25'b1111111110111011110010011;
    rom[2566] = 25'b1111111110011011001011110;
    rom[2567] = 25'b1111111101111010110101001;
    rom[2568] = 25'b1111111101011010101111010;
    rom[2569] = 25'b1111111100111010111010100;
    rom[2570] = 25'b1111111100011011010111101;
    rom[2571] = 25'b1111111011111100000111010;
    rom[2572] = 25'b1111111011011101001001110;
    rom[2573] = 25'b1111111010111110011111110;
    rom[2574] = 25'b1111111010100000001001111;
    rom[2575] = 25'b1111111010000010001000100;
    rom[2576] = 25'b1111111001100100011100010;
    rom[2577] = 25'b1111111001000111000101101;
    rom[2578] = 25'b1111111000101010000101001;
    rom[2579] = 25'b1111111000001101011011011;
    rom[2580] = 25'b1111110111110001001000100;
    rom[2581] = 25'b1111110111010101001101010;
    rom[2582] = 25'b1111110110111001101010001;
    rom[2583] = 25'b1111110110011110011111011;
    rom[2584] = 25'b1111110110000011101101100;
    rom[2585] = 25'b1111110101101001010100111;
    rom[2586] = 25'b1111110101001111010110001;
    rom[2587] = 25'b1111110100110101110001011;
    rom[2588] = 25'b1111110100011100100111010;
    rom[2589] = 25'b1111110100000011110111111;
    rom[2590] = 25'b1111110011101011100011111;
    rom[2591] = 25'b1111110011010011101011100;
    rom[2592] = 25'b1111110010111100001111000;
    rom[2593] = 25'b1111110010100101001110111;
    rom[2594] = 25'b1111110010001110101011010;
    rom[2595] = 25'b1111110001111000100100101;
    rom[2596] = 25'b1111110001100010111011001;
    rom[2597] = 25'b1111110001001101101111010;
    rom[2598] = 25'b1111110000111001000001000;
    rom[2599] = 25'b1111110000100100110000111;
    rom[2600] = 25'b1111110000010000111110111;
    rom[2601] = 25'b1111101111111101101011100;
    rom[2602] = 25'b1111101111101010110110111;
    rom[2603] = 25'b1111101111011000100001001;
    rom[2604] = 25'b1111101111000110101010011;
    rom[2605] = 25'b1111101110110101010011010;
    rom[2606] = 25'b1111101110100100011011011;
    rom[2607] = 25'b1111101110010100000011010;
    rom[2608] = 25'b1111101110000100001011000;
    rom[2609] = 25'b1111101101110100110010101;
    rom[2610] = 25'b1111101101100101111010100;
    rom[2611] = 25'b1111101101010111100010011;
    rom[2612] = 25'b1111101101001001101010110;
    rom[2613] = 25'b1111101100111100010011011;
    rom[2614] = 25'b1111101100101111011100100;
    rom[2615] = 25'b1111101100100011000110010;
    rom[2616] = 25'b1111101100010111010000101;
    rom[2617] = 25'b1111101100001011111011100;
    rom[2618] = 25'b1111101100000001000111010;
    rom[2619] = 25'b1111101011110110110011101;
    rom[2620] = 25'b1111101011101101000000110;
    rom[2621] = 25'b1111101011100011101110101;
    rom[2622] = 25'b1111101011011010111101010;
    rom[2623] = 25'b1111101011010010101100100;
    rom[2624] = 25'b1111101011001010111100100;
    rom[2625] = 25'b1111101011000011101101001;
    rom[2626] = 25'b1111101010111100111110010;
    rom[2627] = 25'b1111101010110110110000000;
    rom[2628] = 25'b1111101010110001000010001;
    rom[2629] = 25'b1111101010101011110100101;
    rom[2630] = 25'b1111101010100111000111010;
    rom[2631] = 25'b1111101010100010111010001;
    rom[2632] = 25'b1111101010011111001101000;
    rom[2633] = 25'b1111101010011011111111111;
    rom[2634] = 25'b1111101010011001010010011;
    rom[2635] = 25'b1111101010010111000100101;
    rom[2636] = 25'b1111101010010101010110010;
    rom[2637] = 25'b1111101010010100000111001;
    rom[2638] = 25'b1111101010010011010111001;
    rom[2639] = 25'b1111101010010011000110001;
    rom[2640] = 25'b1111101010010011010011111;
    rom[2641] = 25'b1111101010010100000000000;
    rom[2642] = 25'b1111101010010101001010101;
    rom[2643] = 25'b1111101010010110110011001;
    rom[2644] = 25'b1111101010011000111001101;
    rom[2645] = 25'b1111101010011011011101110;
    rom[2646] = 25'b1111101010011110011111010;
    rom[2647] = 25'b1111101010100001111101111;
    rom[2648] = 25'b1111101010100101111001010;
    rom[2649] = 25'b1111101010101010010001010;
    rom[2650] = 25'b1111101010101111000101100;
    rom[2651] = 25'b1111101010110100010101110;
    rom[2652] = 25'b1111101010111010000001110;
    rom[2653] = 25'b1111101011000000001001000;
    rom[2654] = 25'b1111101011000110101011100;
    rom[2655] = 25'b1111101011001101101000101;
    rom[2656] = 25'b1111101011010101000000010;
    rom[2657] = 25'b1111101011011100110010000;
    rom[2658] = 25'b1111101011100100111101011;
    rom[2659] = 25'b1111101011101101100010010;
    rom[2660] = 25'b1111101011110110100000001;
    rom[2661] = 25'b1111101011111111110110110;
    rom[2662] = 25'b1111101100001001100101101;
    rom[2663] = 25'b1111101100010011101100100;
    rom[2664] = 25'b1111101100011110001011000;
    rom[2665] = 25'b1111101100101001000000101;
    rom[2666] = 25'b1111101100110100001101000;
    rom[2667] = 25'b1111101100111111101111110;
    rom[2668] = 25'b1111101101001011101000100;
    rom[2669] = 25'b1111101101010111110111000;
    rom[2670] = 25'b1111101101100100011010100;
    rom[2671] = 25'b1111101101110001010010111;
    rom[2672] = 25'b1111101101111110011111101;
    rom[2673] = 25'b1111101110001100000000010;
    rom[2674] = 25'b1111101110011001110100010;
    rom[2675] = 25'b1111101110100111111011100;
    rom[2676] = 25'b1111101110110110010101010;
    rom[2677] = 25'b1111101111000101000001010;
    rom[2678] = 25'b1111101111010011111111000;
    rom[2679] = 25'b1111101111100011001110000;
    rom[2680] = 25'b1111101111110010101110000;
    rom[2681] = 25'b1111110000000010011110010;
    rom[2682] = 25'b1111110000010010011110100;
    rom[2683] = 25'b1111110000100010101110001;
    rom[2684] = 25'b1111110000110011001100111;
    rom[2685] = 25'b1111110001000011111010010;
    rom[2686] = 25'b1111110001010100110101101;
    rom[2687] = 25'b1111110001100101111110101;
    rom[2688] = 25'b1111110001110111010100111;
    rom[2689] = 25'b1111110010001000110111110;
    rom[2690] = 25'b1111110010011010100110111;
    rom[2691] = 25'b1111110010101100100001110;
    rom[2692] = 25'b1111110010111110100111111;
    rom[2693] = 25'b1111110011010000111000111;
    rom[2694] = 25'b1111110011100011010100001;
    rom[2695] = 25'b1111110011110101111001011;
    rom[2696] = 25'b1111110100001000100111111;
    rom[2697] = 25'b1111110100011011011111011;
    rom[2698] = 25'b1111110100101110011111001;
    rom[2699] = 25'b1111110101000001100111000;
    rom[2700] = 25'b1111110101010100110110011;
    rom[2701] = 25'b1111110101101000001100101;
    rom[2702] = 25'b1111110101111011101001101;
    rom[2703] = 25'b1111110110001111001100100;
    rom[2704] = 25'b1111110110100010110101000;
    rom[2705] = 25'b1111110110110110100010110;
    rom[2706] = 25'b1111110111001010010101000;
    rom[2707] = 25'b1111110111011110001011100;
    rom[2708] = 25'b1111110111110010000101101;
    rom[2709] = 25'b1111111000000110000011001;
    rom[2710] = 25'b1111111000011010000011011;
    rom[2711] = 25'b1111111000101110000101111;
    rom[2712] = 25'b1111111001000010001010011;
    rom[2713] = 25'b1111111001010110010000001;
    rom[2714] = 25'b1111111001101010010111000;
    rom[2715] = 25'b1111111001111110011110011;
    rom[2716] = 25'b1111111010010010100101101;
    rom[2717] = 25'b1111111010100110101100101;
    rom[2718] = 25'b1111111010111010110010110;
    rom[2719] = 25'b1111111011001110110111101;
    rom[2720] = 25'b1111111011100010111010110;
    rom[2721] = 25'b1111111011110110111011111;
    rom[2722] = 25'b1111111100001010111010011;
    rom[2723] = 25'b1111111100011110110101110;
    rom[2724] = 25'b1111111100110010101101111;
    rom[2725] = 25'b1111111101000110100010001;
    rom[2726] = 25'b1111111101011010010010001;
    rom[2727] = 25'b1111111101101101111101011;
    rom[2728] = 25'b1111111110000001100011110;
    rom[2729] = 25'b1111111110010101000100100;
    rom[2730] = 25'b1111111110101000011111100;
    rom[2731] = 25'b1111111110111011110100010;
    rom[2732] = 25'b1111111111001111000010010;
    rom[2733] = 25'b1111111111100010001001010;
    rom[2734] = 25'b1111111111110101001000111;
    rom[2735] = 25'b0000000000001000000000101;
    rom[2736] = 25'b0000000000011010110000011;
    rom[2737] = 25'b0000000000101101010111101;
    rom[2738] = 25'b0000000000111111110110000;
    rom[2739] = 25'b0000000001010010001011010;
    rom[2740] = 25'b0000000001100100010110111;
    rom[2741] = 25'b0000000001110110011000101;
    rom[2742] = 25'b0000000010001000010000000;
    rom[2743] = 25'b0000000010011001111101000;
    rom[2744] = 25'b0000000010101011011111000;
    rom[2745] = 25'b0000000010111100110101111;
    rom[2746] = 25'b0000000011001110000001010;
    rom[2747] = 25'b0000000011011111000000110;
    rom[2748] = 25'b0000000011101111110100010;
    rom[2749] = 25'b0000000100000000011011001;
    rom[2750] = 25'b0000000100010000110101100;
    rom[2751] = 25'b0000000100100001000010111;
    rom[2752] = 25'b0000000100110001000011000;
    rom[2753] = 25'b0000000101000000110101100;
    rom[2754] = 25'b0000000101010000011010010;
    rom[2755] = 25'b0000000101011111110001001;
    rom[2756] = 25'b0000000101101110111001101;
    rom[2757] = 25'b0000000101111101110011101;
    rom[2758] = 25'b0000000110001100011110110;
    rom[2759] = 25'b0000000110011010111011000;
    rom[2760] = 25'b0000000110101001001000000;
    rom[2761] = 25'b0000000110110111000101101;
    rom[2762] = 25'b0000000111000100110011100;
    rom[2763] = 25'b0000000111010010010001101;
    rom[2764] = 25'b0000000111011111011111110;
    rom[2765] = 25'b0000000111101100011101110;
    rom[2766] = 25'b0000000111111001001011001;
    rom[2767] = 25'b0000001000000101101000000;
    rom[2768] = 25'b0000001000010001110100010;
    rom[2769] = 25'b0000001000011101101111100;
    rom[2770] = 25'b0000001000101001011001110;
    rom[2771] = 25'b0000001000110100110010111;
    rom[2772] = 25'b0000001000111111111010011;
    rom[2773] = 25'b0000001001001010110000110;
    rom[2774] = 25'b0000001001010101010101011;
    rom[2775] = 25'b0000001001011111101000010;
    rom[2776] = 25'b0000001001101001101001011;
    rom[2777] = 25'b0000001001110011011000100;
    rom[2778] = 25'b0000001001111100110101101;
    rom[2779] = 25'b0000001010000110000000101;
    rom[2780] = 25'b0000001010001110111001100;
    rom[2781] = 25'b0000001010010111100000001;
    rom[2782] = 25'b0000001010011111110100010;
    rom[2783] = 25'b0000001010100111110110001;
    rom[2784] = 25'b0000001010101111100101011;
    rom[2785] = 25'b0000001010110111000010001;
    rom[2786] = 25'b0000001010111110001100011;
    rom[2787] = 25'b0000001011000101000100001;
    rom[2788] = 25'b0000001011001011101001000;
    rom[2789] = 25'b0000001011010001111011100;
    rom[2790] = 25'b0000001011010111111011001;
    rom[2791] = 25'b0000001011011101101000001;
    rom[2792] = 25'b0000001011100011000010100;
    rom[2793] = 25'b0000001011101000001010001;
    rom[2794] = 25'b0000001011101100111111001;
    rom[2795] = 25'b0000001011110001100001100;
    rom[2796] = 25'b0000001011110101110001011;
    rom[2797] = 25'b0000001011111001101110011;
    rom[2798] = 25'b0000001011111101011001000;
    rom[2799] = 25'b0000001100000000110001001;
    rom[2800] = 25'b0000001100000011110110110;
    rom[2801] = 25'b0000001100000110101001111;
    rom[2802] = 25'b0000001100001001001010110;
    rom[2803] = 25'b0000001100001011011001011;
    rom[2804] = 25'b0000001100001101010101101;
    rom[2805] = 25'b0000001100001110111111111;
    rom[2806] = 25'b0000001100010000011000000;
    rom[2807] = 25'b0000001100010001011110001;
    rom[2808] = 25'b0000001100010010010010100;
    rom[2809] = 25'b0000001100010010110101000;
    rom[2810] = 25'b0000001100010011000101111;
    rom[2811] = 25'b0000001100010011000101010;
    rom[2812] = 25'b0000001100010010110011001;
    rom[2813] = 25'b0000001100010010001111110;
    rom[2814] = 25'b0000001100010001011011001;
    rom[2815] = 25'b0000001100010000010101100;
    rom[2816] = 25'b0000001100001110111111000;
    rom[2817] = 25'b0000001100001101010111110;
    rom[2818] = 25'b0000001100001011011111110;
    rom[2819] = 25'b0000001100001001010111011;
    rom[2820] = 25'b0000001100000110111110101;
    rom[2821] = 25'b0000001100000100010101111;
    rom[2822] = 25'b0000001100000001011101000;
    rom[2823] = 25'b0000001011111110010100011;
    rom[2824] = 25'b0000001011111010111100001;
    rom[2825] = 25'b0000001011110111010100011;
    rom[2826] = 25'b0000001011110011011101100;
    rom[2827] = 25'b0000001011101111010111011;
    rom[2828] = 25'b0000001011101011000010011;
    rom[2829] = 25'b0000001011100110011110111;
    rom[2830] = 25'b0000001011100001101100110;
    rom[2831] = 25'b0000001011011100101100011;
    rom[2832] = 25'b0000001011010111011101110;
    rom[2833] = 25'b0000001011010010000001011;
    rom[2834] = 25'b0000001011001100010111100;
    rom[2835] = 25'b0000001011000110100000000;
    rom[2836] = 25'b0000001011000000011011011;
    rom[2837] = 25'b0000001010111010001001110;
    rom[2838] = 25'b0000001010110011101011011;
    rom[2839] = 25'b0000001010101101000000011;
    rom[2840] = 25'b0000001010100110001001010;
    rom[2841] = 25'b0000001010011111000101111;
    rom[2842] = 25'b0000001010010111110110110;
    rom[2843] = 25'b0000001010010000011100000;
    rom[2844] = 25'b0000001010001000110110000;
    rom[2845] = 25'b0000001010000001000100111;
    rom[2846] = 25'b0000001001111001001000110;
    rom[2847] = 25'b0000001001110001000010010;
    rom[2848] = 25'b0000001001101000110001011;
    rom[2849] = 25'b0000001001100000010110011;
    rom[2850] = 25'b0000001001010111110001100;
    rom[2851] = 25'b0000001001001111000011000;
    rom[2852] = 25'b0000001001000110001011011;
    rom[2853] = 25'b0000001000111101001010100;
    rom[2854] = 25'b0000001000110100000001000;
    rom[2855] = 25'b0000001000101010101110110;
    rom[2856] = 25'b0000001000100001010100011;
    rom[2857] = 25'b0000001000010111110010000;
    rom[2858] = 25'b0000001000001110000111111;
    rom[2859] = 25'b0000001000000100010110011;
    rom[2860] = 25'b0000000111111010011101101;
    rom[2861] = 25'b0000000111110000011110000;
    rom[2862] = 25'b0000000111100110010111101;
    rom[2863] = 25'b0000000111011100001010111;
    rom[2864] = 25'b0000000111010001111000000;
    rom[2865] = 25'b0000000111000111011111010;
    rom[2866] = 25'b0000000110111101000001001;
    rom[2867] = 25'b0000000110110010011101100;
    rom[2868] = 25'b0000000110100111110100111;
    rom[2869] = 25'b0000000110011101000111100;
    rom[2870] = 25'b0000000110010010010101110;
    rom[2871] = 25'b0000000110000111011111110;
    rom[2872] = 25'b0000000101111100100101110;
    rom[2873] = 25'b0000000101110001101000001;
    rom[2874] = 25'b0000000101100110100111000;
    rom[2875] = 25'b0000000101011011100010111;
    rom[2876] = 25'b0000000101010000011011110;
    rom[2877] = 25'b0000000101000101010010001;
    rom[2878] = 25'b0000000100111010000110010;
    rom[2879] = 25'b0000000100101110111000001;
    rom[2880] = 25'b0000000100100011101000011;
    rom[2881] = 25'b0000000100011000010111000;
    rom[2882] = 25'b0000000100001101000100011;
    rom[2883] = 25'b0000000100000001110000110;
    rom[2884] = 25'b0000000011110110011100010;
    rom[2885] = 25'b0000000011101011000111011;
    rom[2886] = 25'b0000000011011111110010010;
    rom[2887] = 25'b0000000011010100011101001;
    rom[2888] = 25'b0000000011001001001000010;
    rom[2889] = 25'b0000000010111101110100000;
    rom[2890] = 25'b0000000010110010100000011;
    rom[2891] = 25'b0000000010100111001101111;
    rom[2892] = 25'b0000000010011011111100101;
    rom[2893] = 25'b0000000010010000101100110;
    rom[2894] = 25'b0000000010000101011110111;
    rom[2895] = 25'b0000000001111010010010110;
    rom[2896] = 25'b0000000001101111001001000;
    rom[2897] = 25'b0000000001100100000001101;
    rom[2898] = 25'b0000000001011000111101000;
    rom[2899] = 25'b0000000001001101111011010;
    rom[2900] = 25'b0000000001000010111100101;
    rom[2901] = 25'b0000000000111000000001011;
    rom[2902] = 25'b0000000000101101001001111;
    rom[2903] = 25'b0000000000100010010110000;
    rom[2904] = 25'b0000000000010111100110010;
    rom[2905] = 25'b0000000000001100111010101;
    rom[2906] = 25'b0000000000000010010011101;
    rom[2907] = 25'b1111111111110111110001001;
    rom[2908] = 25'b1111111111101101010011101;
    rom[2909] = 25'b1111111111100010111011000;
    rom[2910] = 25'b1111111111011000100111110;
    rom[2911] = 25'b1111111111001110011001111;
    rom[2912] = 25'b1111111111000100010001110;
    rom[2913] = 25'b1111111110111010001111011;
    rom[2914] = 25'b1111111110110000010011000;
    rom[2915] = 25'b1111111110100110011100111;
    rom[2916] = 25'b1111111110011100101101001;
    rom[2917] = 25'b1111111110010011000011111;
    rom[2918] = 25'b1111111110001001100001011;
    rom[2919] = 25'b1111111110000000000101110;
    rom[2920] = 25'b1111111101110110110001001;
    rom[2921] = 25'b1111111101101101100011110;
    rom[2922] = 25'b1111111101100100011101110;
    rom[2923] = 25'b1111111101011011011111010;
    rom[2924] = 25'b1111111101010010101000011;
    rom[2925] = 25'b1111111101001001111001011;
    rom[2926] = 25'b1111111101000001010010011;
    rom[2927] = 25'b1111111100111000110011011;
    rom[2928] = 25'b1111111100110000011100101;
    rom[2929] = 25'b1111111100101000001110010;
    rom[2930] = 25'b1111111100100000001000010;
    rom[2931] = 25'b1111111100011000001011000;
    rom[2932] = 25'b1111111100010000010110010;
    rom[2933] = 25'b1111111100001000101010101;
    rom[2934] = 25'b1111111100000001000111110;
    rom[2935] = 25'b1111111011111001101101111;
    rom[2936] = 25'b1111111011110010011101011;
    rom[2937] = 25'b1111111011101011010110000;
    rom[2938] = 25'b1111111011100100010111111;
    rom[2939] = 25'b1111111011011101100011011;
    rom[2940] = 25'b1111111011010110111000010;
    rom[2941] = 25'b1111111011010000010110111;
    rom[2942] = 25'b1111111011001001111111001;
    rom[2943] = 25'b1111111011000011110001001;
    rom[2944] = 25'b1111111010111101101100111;
    rom[2945] = 25'b1111111010110111110010101;
    rom[2946] = 25'b1111111010110010000010011;
    rom[2947] = 25'b1111111010101100011100001;
    rom[2948] = 25'b1111111010100111000000000;
    rom[2949] = 25'b1111111010100001101101111;
    rom[2950] = 25'b1111111010011100100110000;
    rom[2951] = 25'b1111111010010111101000011;
    rom[2952] = 25'b1111111010010010110100111;
    rom[2953] = 25'b1111111010001110001011111;
    rom[2954] = 25'b1111111010001001101101001;
    rom[2955] = 25'b1111111010000101011000101;
    rom[2956] = 25'b1111111010000001001110101;
    rom[2957] = 25'b1111111001111101001111000;
    rom[2958] = 25'b1111111001111001011001111;
    rom[2959] = 25'b1111111001110101101111000;
    rom[2960] = 25'b1111111001110010001110101;
    rom[2961] = 25'b1111111001101110111000110;
    rom[2962] = 25'b1111111001101011101101011;
    rom[2963] = 25'b1111111001101000101100010;
    rom[2964] = 25'b1111111001100101110101110;
    rom[2965] = 25'b1111111001100011001001101;
    rom[2966] = 25'b1111111001100000100111111;
    rom[2967] = 25'b1111111001011110010000100;
    rom[2968] = 25'b1111111001011100000011100;
    rom[2969] = 25'b1111111001011010000000111;
    rom[2970] = 25'b1111111001011000001000101;
    rom[2971] = 25'b1111111001010110011010101;
    rom[2972] = 25'b1111111001010100110110111;
    rom[2973] = 25'b1111111001010011011101100;
    rom[2974] = 25'b1111111001010010001110001;
    rom[2975] = 25'b1111111001010001001001000;
    rom[2976] = 25'b1111111001010000001101111;
    rom[2977] = 25'b1111111001001111011100111;
    rom[2978] = 25'b1111111001001110110101110;
    rom[2979] = 25'b1111111001001110011000101;
    rom[2980] = 25'b1111111001001110000101011;
    rom[2981] = 25'b1111111001001101111100000;
    rom[2982] = 25'b1111111001001101111100010;
    rom[2983] = 25'b1111111001001110000110010;
    rom[2984] = 25'b1111111001001110011001110;
    rom[2985] = 25'b1111111001001110110110110;
    rom[2986] = 25'b1111111001001111011101010;
    rom[2987] = 25'b1111111001010000001101010;
    rom[2988] = 25'b1111111001010001000110011;
    rom[2989] = 25'b1111111001010010001000110;
    rom[2990] = 25'b1111111001010011010100001;
    rom[2991] = 25'b1111111001010100101000101;
    rom[2992] = 25'b1111111001010110000110000;
    rom[2993] = 25'b1111111001010111101100010;
    rom[2994] = 25'b1111111001011001011011001;
    rom[2995] = 25'b1111111001011011010010110;
    rom[2996] = 25'b1111111001011101010010111;
    rom[2997] = 25'b1111111001011111011011011;
    rom[2998] = 25'b1111111001100001101100001;
    rom[2999] = 25'b1111111001100100000101001;
    rom[3000] = 25'b1111111001100110100110001;
    rom[3001] = 25'b1111111001101001001111010;
    rom[3002] = 25'b1111111001101100000000001;
    rom[3003] = 25'b1111111001101110111000110;
    rom[3004] = 25'b1111111001110001111001000;
    rom[3005] = 25'b1111111001110101000000101;
    rom[3006] = 25'b1111111001111000001111111;
    rom[3007] = 25'b1111111001111011100110001;
    rom[3008] = 25'b1111111001111111000011101;
    rom[3009] = 25'b1111111010000010101000001;
    rom[3010] = 25'b1111111010000110010011011;
    rom[3011] = 25'b1111111010001010000101011;
    rom[3012] = 25'b1111111010001101111110000;
    rom[3013] = 25'b1111111010010001111101000;
    rom[3014] = 25'b1111111010010110000010011;
    rom[3015] = 25'b1111111010011010001101111;
    rom[3016] = 25'b1111111010011110011111100;
    rom[3017] = 25'b1111111010100010110111000;
    rom[3018] = 25'b1111111010100111010100010;
    rom[3019] = 25'b1111111010101011110111001;
    rom[3020] = 25'b1111111010110000011111100;
    rom[3021] = 25'b1111111010110101001101010;
    rom[3022] = 25'b1111111010111010000000001;
    rom[3023] = 25'b1111111010111110111000000;
    rom[3024] = 25'b1111111011000011110100110;
    rom[3025] = 25'b1111111011001000110110011;
    rom[3026] = 25'b1111111011001101111100101;
    rom[3027] = 25'b1111111011010011000111010;
    rom[3028] = 25'b1111111011011000010110001;
    rom[3029] = 25'b1111111011011101101001001;
    rom[3030] = 25'b1111111011100011000000010;
    rom[3031] = 25'b1111111011101000011011010;
    rom[3032] = 25'b1111111011101101111001111;
    rom[3033] = 25'b1111111011110011011100000;
    rom[3034] = 25'b1111111011111001000001110;
    rom[3035] = 25'b1111111011111110101010101;
    rom[3036] = 25'b1111111100000100010110101;
    rom[3037] = 25'b1111111100001010000101100;
    rom[3038] = 25'b1111111100001111110111001;
    rom[3039] = 25'b1111111100010101101011101;
    rom[3040] = 25'b1111111100011011100010100;
    rom[3041] = 25'b1111111100100001011011110;
    rom[3042] = 25'b1111111100100111010111010;
    rom[3043] = 25'b1111111100101101010100101;
    rom[3044] = 25'b1111111100110011010100000;
    rom[3045] = 25'b1111111100111001010101010;
    rom[3046] = 25'b1111111100111111011000000;
    rom[3047] = 25'b1111111101000101011100010;
    rom[3048] = 25'b1111111101001011100001110;
    rom[3049] = 25'b1111111101010001101000100;
    rom[3050] = 25'b1111111101010111110000010;
    rom[3051] = 25'b1111111101011101111000110;
    rom[3052] = 25'b1111111101100100000010001;
    rom[3053] = 25'b1111111101101010001100000;
    rom[3054] = 25'b1111111101110000010110011;
    rom[3055] = 25'b1111111101110110100001000;
    rom[3056] = 25'b1111111101111100101011111;
    rom[3057] = 25'b1111111110000010110110101;
    rom[3058] = 25'b1111111110001001000001010;
    rom[3059] = 25'b1111111110001111001011110;
    rom[3060] = 25'b1111111110010101010101110;
    rom[3061] = 25'b1111111110011011011111011;
    rom[3062] = 25'b1111111110100001101000001;
    rom[3063] = 25'b1111111110100111110000010;
    rom[3064] = 25'b1111111110101101110111010;
    rom[3065] = 25'b1111111110110011111101011;
    rom[3066] = 25'b1111111110111010000010010;
    rom[3067] = 25'b1111111111000000000101110;
    rom[3068] = 25'b1111111111000110000111110;
    rom[3069] = 25'b1111111111001100001000011;
    rom[3070] = 25'b1111111111010010000111001;
    rom[3071] = 25'b1111111111011000000100001;
    rom[3072] = 25'b1111111111011101111111001;
    rom[3073] = 25'b1111111111100011111000010;
    rom[3074] = 25'b1111111111101001101111000;
    rom[3075] = 25'b1111111111101111100011100;
    rom[3076] = 25'b1111111111110101010101101;
    rom[3077] = 25'b1111111111111011000101010;
    rom[3078] = 25'b0000000000000000110010001;
    rom[3079] = 25'b0000000000000110011100010;
    rom[3080] = 25'b0000000000001100000011101;
    rom[3081] = 25'b0000000000010001101000000;
    rom[3082] = 25'b0000000000010111001001011;
    rom[3083] = 25'b0000000000011100100111101;
    rom[3084] = 25'b0000000000100010000010100;
    rom[3085] = 25'b0000000000100111011010001;
    rom[3086] = 25'b0000000000101100101110010;
    rom[3087] = 25'b0000000000110001111110111;
    rom[3088] = 25'b0000000000110111001011110;
    rom[3089] = 25'b0000000000111100010101000;
    rom[3090] = 25'b0000000001000001011010011;
    rom[3091] = 25'b0000000001000110011011110;
    rom[3092] = 25'b0000000001001011011001010;
    rom[3093] = 25'b0000000001010000010010101;
    rom[3094] = 25'b0000000001010101001000000;
    rom[3095] = 25'b0000000001011001111001001;
    rom[3096] = 25'b0000000001011110100101110;
    rom[3097] = 25'b0000000001100011001110001;
    rom[3098] = 25'b0000000001100111110010000;
    rom[3099] = 25'b0000000001101100010001011;
    rom[3100] = 25'b0000000001110000101100001;
    rom[3101] = 25'b0000000001110101000010010;
    rom[3102] = 25'b0000000001111001010011101;
    rom[3103] = 25'b0000000001111101100000010;
    rom[3104] = 25'b0000000010000001101000001;
    rom[3105] = 25'b0000000010000101101011000;
    rom[3106] = 25'b0000000010001001101001000;
    rom[3107] = 25'b0000000010001101100001111;
    rom[3108] = 25'b0000000010010001010101110;
    rom[3109] = 25'b0000000010010101000100101;
    rom[3110] = 25'b0000000010011000101110010;
    rom[3111] = 25'b0000000010011100010010110;
    rom[3112] = 25'b0000000010011111110010000;
    rom[3113] = 25'b0000000010100011001011111;
    rom[3114] = 25'b0000000010100110100000100;
    rom[3115] = 25'b0000000010101001101111111;
    rom[3116] = 25'b0000000010101100111001110;
    rom[3117] = 25'b0000000010101111111110010;
    rom[3118] = 25'b0000000010110010111101011;
    rom[3119] = 25'b0000000010110101110110111;
    rom[3120] = 25'b0000000010111000101011001;
    rom[3121] = 25'b0000000010111011011001110;
    rom[3122] = 25'b0000000010111110000010110;
    rom[3123] = 25'b0000000011000000100110011;
    rom[3124] = 25'b0000000011000011000100010;
    rom[3125] = 25'b0000000011000101011100111;
    rom[3126] = 25'b0000000011000111101111101;
    rom[3127] = 25'b0000000011001001111100111;
    rom[3128] = 25'b0000000011001100000100100;
    rom[3129] = 25'b0000000011001110000110011;
    rom[3130] = 25'b0000000011010000000010111;
    rom[3131] = 25'b0000000011010001111001101;
    rom[3132] = 25'b0000000011010011101010110;
    rom[3133] = 25'b0000000011010101010110011;
    rom[3134] = 25'b0000000011010110111100011;
    rom[3135] = 25'b0000000011011000011100101;
    rom[3136] = 25'b0000000011011001110111011;
    rom[3137] = 25'b0000000011011011001100101;
    rom[3138] = 25'b0000000011011100011100010;
    rom[3139] = 25'b0000000011011101100110010;
    rom[3140] = 25'b0000000011011110101010110;
    rom[3141] = 25'b0000000011011111101001110;
    rom[3142] = 25'b0000000011100000100011010;
    rom[3143] = 25'b0000000011100001010111010;
    rom[3144] = 25'b0000000011100010000101111;
    rom[3145] = 25'b0000000011100010101111000;
    rom[3146] = 25'b0000000011100011010010111;
    rom[3147] = 25'b0000000011100011110001001;
    rom[3148] = 25'b0000000011100100001010001;
    rom[3149] = 25'b0000000011100100011101111;
    rom[3150] = 25'b0000000011100100101100010;
    rom[3151] = 25'b0000000011100100110101100;
    rom[3152] = 25'b0000000011100100111001100;
    rom[3153] = 25'b0000000011100100111000011;
    rom[3154] = 25'b0000000011100100110010000;
    rom[3155] = 25'b0000000011100100100110101;
    rom[3156] = 25'b0000000011100100010110010;
    rom[3157] = 25'b0000000011100100000000110;
    rom[3158] = 25'b0000000011100011100110011;
    rom[3159] = 25'b0000000011100011000111001;
    rom[3160] = 25'b0000000011100010100010111;
    rom[3161] = 25'b0000000011100001111010000;
    rom[3162] = 25'b0000000011100001001100010;
    rom[3163] = 25'b0000000011100000011001111;
    rom[3164] = 25'b0000000011011111100010111;
    rom[3165] = 25'b0000000011011110100111010;
    rom[3166] = 25'b0000000011011101100111001;
    rom[3167] = 25'b0000000011011100100010100;
    rom[3168] = 25'b0000000011011011011001011;
    rom[3169] = 25'b0000000011011010001100000;
    rom[3170] = 25'b0000000011011000111010010;
    rom[3171] = 25'b0000000011010111100100011;
    rom[3172] = 25'b0000000011010110001010010;
    rom[3173] = 25'b0000000011010100101100000;
    rom[3174] = 25'b0000000011010011001001110;
    rom[3175] = 25'b0000000011010001100011100;
    rom[3176] = 25'b0000000011001111111001011;
    rom[3177] = 25'b0000000011001110001011011;
    rom[3178] = 25'b0000000011001100011001101;
    rom[3179] = 25'b0000000011001010100100010;
    rom[3180] = 25'b0000000011001000101011001;
    rom[3181] = 25'b0000000011000110101110100;
    rom[3182] = 25'b0000000011000100101110011;
    rom[3183] = 25'b0000000011000010101010111;
    rom[3184] = 25'b0000000011000000100100000;
    rom[3185] = 25'b0000000010111110011001111;
    rom[3186] = 25'b0000000010111100001100011;
    rom[3187] = 25'b0000000010111001111100000;
    rom[3188] = 25'b0000000010110111101000100;
    rom[3189] = 25'b0000000010110101010010000;
    rom[3190] = 25'b0000000010110010111000101;
    rom[3191] = 25'b0000000010110000011100100;
    rom[3192] = 25'b0000000010101101111101101;
    rom[3193] = 25'b0000000010101011011100000;
    rom[3194] = 25'b0000000010101000110111111;
    rom[3195] = 25'b0000000010100110010001010;
    rom[3196] = 25'b0000000010100011101000001;
    rom[3197] = 25'b0000000010100000111100110;
    rom[3198] = 25'b0000000010011110001111000;
    rom[3199] = 25'b0000000010011011011111010;
    rom[3200] = 25'b0000000010011000101101010;
    rom[3201] = 25'b0000000010010101111001010;
    rom[3202] = 25'b0000000010010011000011011;
    rom[3203] = 25'b0000000010010000001011100;
    rom[3204] = 25'b0000000010001101010001111;
    rom[3205] = 25'b0000000010001010010110101;
    rom[3206] = 25'b0000000010000111011001110;
    rom[3207] = 25'b0000000010000100011011010;
    rom[3208] = 25'b0000000010000001011011011;
    rom[3209] = 25'b0000000001111110011010000;
    rom[3210] = 25'b0000000001111011010111011;
    rom[3211] = 25'b0000000001111000010011100;
    rom[3212] = 25'b0000000001110101001110100;
    rom[3213] = 25'b0000000001110010001000100;
    rom[3214] = 25'b0000000001101111000001011;
    rom[3215] = 25'b0000000001101011111001011;
    rom[3216] = 25'b0000000001101000110000101;
    rom[3217] = 25'b0000000001100101100111001;
    rom[3218] = 25'b0000000001100010011100110;
    rom[3219] = 25'b0000000001011111010010000;
    rom[3220] = 25'b0000000001011100000110101;
    rom[3221] = 25'b0000000001011000111010110;
    rom[3222] = 25'b0000000001010101101110100;
    rom[3223] = 25'b0000000001010010100010001;
    rom[3224] = 25'b0000000001001111010101011;
    rom[3225] = 25'b0000000001001100001000100;
    rom[3226] = 25'b0000000001001000111011100;
    rom[3227] = 25'b0000000001000101101110101;
    rom[3228] = 25'b0000000001000010100001110;
    rom[3229] = 25'b0000000000111111010101001;
    rom[3230] = 25'b0000000000111100001000101;
    rom[3231] = 25'b0000000000111000111100011;
    rom[3232] = 25'b0000000000110101110000100;
    rom[3233] = 25'b0000000000110010100101001;
    rom[3234] = 25'b0000000000101111011010010;
    rom[3235] = 25'b0000000000101100001111111;
    rom[3236] = 25'b0000000000101001000110001;
    rom[3237] = 25'b0000000000100101111101001;
    rom[3238] = 25'b0000000000100010110100111;
    rom[3239] = 25'b0000000000011111101101100;
    rom[3240] = 25'b0000000000011100100110111;
    rom[3241] = 25'b0000000000011001100001010;
    rom[3242] = 25'b0000000000010110011100110;
    rom[3243] = 25'b0000000000010011011001010;
    rom[3244] = 25'b0000000000010000010111000;
    rom[3245] = 25'b0000000000001101010101110;
    rom[3246] = 25'b0000000000001010010101111;
    rom[3247] = 25'b0000000000000111010111011;
    rom[3248] = 25'b0000000000000100011010010;
    rom[3249] = 25'b0000000000000001011110100;
    rom[3250] = 25'b1111111111111110100100010;
    rom[3251] = 25'b1111111111111011101011100;
    rom[3252] = 25'b1111111111111000110100011;
    rom[3253] = 25'b1111111111110101111111000;
    rom[3254] = 25'b1111111111110011001011001;
    rom[3255] = 25'b1111111111110000011001001;
    rom[3256] = 25'b1111111111101101101001000;
    rom[3257] = 25'b1111111111101010111010100;
    rom[3258] = 25'b1111111111101000001110001;
    rom[3259] = 25'b1111111111100101100011100;
    rom[3260] = 25'b1111111111100010111011000;
    rom[3261] = 25'b1111111111100000010100011;
    rom[3262] = 25'b1111111111011101110000000;
    rom[3263] = 25'b1111111111011011001101101;
    rom[3264] = 25'b1111111111011000101101011;
    rom[3265] = 25'b1111111111010110001111011;
    rom[3266] = 25'b1111111111010011110011101;
    rom[3267] = 25'b1111111111010001011010010;
    rom[3268] = 25'b1111111111001111000011000;
    rom[3269] = 25'b1111111111001100101110001;
    rom[3270] = 25'b1111111111001010011011101;
    rom[3271] = 25'b1111111111001000001011101;
    rom[3272] = 25'b1111111111000101111110000;
    rom[3273] = 25'b1111111111000011110010111;
    rom[3274] = 25'b1111111111000001101010001;
    rom[3275] = 25'b1111111110111111100100000;
    rom[3276] = 25'b1111111110111101100000011;
    rom[3277] = 25'b1111111110111011011111011;
    rom[3278] = 25'b1111111110111001100001001;
    rom[3279] = 25'b1111111110110111100101011;
    rom[3280] = 25'b1111111110110101101100010;
    rom[3281] = 25'b1111111110110011110101110;
    rom[3282] = 25'b1111111110110010000010000;
    rom[3283] = 25'b1111111110110000010001000;
    rom[3284] = 25'b1111111110101110100010110;
    rom[3285] = 25'b1111111110101100110111001;
    rom[3286] = 25'b1111111110101011001110011;
    rom[3287] = 25'b1111111110101001101000010;
    rom[3288] = 25'b1111111110101000000101001;
    rom[3289] = 25'b1111111110100110100100110;
    rom[3290] = 25'b1111111110100101000111001;
    rom[3291] = 25'b1111111110100011101100011;
    rom[3292] = 25'b1111111110100010010100100;
    rom[3293] = 25'b1111111110100000111111011;
    rom[3294] = 25'b1111111110011111101101001;
    rom[3295] = 25'b1111111110011110011101110;
    rom[3296] = 25'b1111111110011101010001001;
    rom[3297] = 25'b1111111110011100000111100;
    rom[3298] = 25'b1111111110011011000000110;
    rom[3299] = 25'b1111111110011001111100111;
    rom[3300] = 25'b1111111110011000111011110;
    rom[3301] = 25'b1111111110010111111101101;
    rom[3302] = 25'b1111111110010111000010010;
    rom[3303] = 25'b1111111110010110001001110;
    rom[3304] = 25'b1111111110010101010100010;
    rom[3305] = 25'b1111111110010100100001100;
    rom[3306] = 25'b1111111110010011110001101;
    rom[3307] = 25'b1111111110010011000100101;
    rom[3308] = 25'b1111111110010010011010011;
    rom[3309] = 25'b1111111110010001110011000;
    rom[3310] = 25'b1111111110010001001110100;
    rom[3311] = 25'b1111111110010000101100110;
    rom[3312] = 25'b1111111110010000001101110;
    rom[3313] = 25'b1111111110001111110001100;
    rom[3314] = 25'b1111111110001111011000001;
    rom[3315] = 25'b1111111110001111000001100;
    rom[3316] = 25'b1111111110001110101101101;
    rom[3317] = 25'b1111111110001110011100100;
    rom[3318] = 25'b1111111110001110001110000;
    rom[3319] = 25'b1111111110001110000010011;
    rom[3320] = 25'b1111111110001101111001001;
    rom[3321] = 25'b1111111110001101110010110;
    rom[3322] = 25'b1111111110001101101111000;
    rom[3323] = 25'b1111111110001101101101110;
    rom[3324] = 25'b1111111110001101101111010;
    rom[3325] = 25'b1111111110001101110011010;
    rom[3326] = 25'b1111111110001101111001110;
    rom[3327] = 25'b1111111110001110000010111;
    rom[3328] = 25'b1111111110001110001110011;
    rom[3329] = 25'b1111111110001110011100100;
    rom[3330] = 25'b1111111110001110101101000;
    rom[3331] = 25'b1111111110001110111111111;
    rom[3332] = 25'b1111111110001111010101001;
    rom[3333] = 25'b1111111110001111101100111;
    rom[3334] = 25'b1111111110010000000111000;
    rom[3335] = 25'b1111111110010000100011010;
    rom[3336] = 25'b1111111110010001000001111;
    rom[3337] = 25'b1111111110010001100010110;
    rom[3338] = 25'b1111111110010010000101111;
    rom[3339] = 25'b1111111110010010101011010;
    rom[3340] = 25'b1111111110010011010010101;
    rom[3341] = 25'b1111111110010011111100010;
    rom[3342] = 25'b1111111110010100100111111;
    rom[3343] = 25'b1111111110010101010101101;
    rom[3344] = 25'b1111111110010110000101011;
    rom[3345] = 25'b1111111110010110110111001;
    rom[3346] = 25'b1111111110010111101010110;
    rom[3347] = 25'b1111111110011000100000100;
    rom[3348] = 25'b1111111110011001010111111;
    rom[3349] = 25'b1111111110011010010001011;
    rom[3350] = 25'b1111111110011011001100100;
    rom[3351] = 25'b1111111110011100001001100;
    rom[3352] = 25'b1111111110011101001000001;
    rom[3353] = 25'b1111111110011110001000100;
    rom[3354] = 25'b1111111110011111001010101;
    rom[3355] = 25'b1111111110100000001110010;
    rom[3356] = 25'b1111111110100001010011101;
    rom[3357] = 25'b1111111110100010011010100;
    rom[3358] = 25'b1111111110100011100010111;
    rom[3359] = 25'b1111111110100100101100101;
    rom[3360] = 25'b1111111110100101111000000;
    rom[3361] = 25'b1111111110100111000100101;
    rom[3362] = 25'b1111111110101000010010101;
    rom[3363] = 25'b1111111110101001100010000;
    rom[3364] = 25'b1111111110101010110010101;
    rom[3365] = 25'b1111111110101100000100100;
    rom[3366] = 25'b1111111110101101010111101;
    rom[3367] = 25'b1111111110101110101011111;
    rom[3368] = 25'b1111111110110000000001001;
    rom[3369] = 25'b1111111110110001010111101;
    rom[3370] = 25'b1111111110110010101111001;
    rom[3371] = 25'b1111111110110100000111100;
    rom[3372] = 25'b1111111110110101100001000;
    rom[3373] = 25'b1111111110110110111011011;
    rom[3374] = 25'b1111111110111000010110100;
    rom[3375] = 25'b1111111110111001110010101;
    rom[3376] = 25'b1111111110111011001111100;
    rom[3377] = 25'b1111111110111100101101000;
    rom[3378] = 25'b1111111110111110001011011;
    rom[3379] = 25'b1111111110111111101010100;
    rom[3380] = 25'b1111111111000001001010001;
    rom[3381] = 25'b1111111111000010101010011;
    rom[3382] = 25'b1111111111000100001011001;
    rom[3383] = 25'b1111111111000101101100100;
    rom[3384] = 25'b1111111111000111001110010;
    rom[3385] = 25'b1111111111001000110000100;
    rom[3386] = 25'b1111111111001010010011010;
    rom[3387] = 25'b1111111111001011110110010;
    rom[3388] = 25'b1111111111001101011001101;
    rom[3389] = 25'b1111111111001110111101010;
    rom[3390] = 25'b1111111111010000100001001;
    rom[3391] = 25'b1111111111010010000101010;
    rom[3392] = 25'b1111111111010011101001011;
    rom[3393] = 25'b1111111111010101001101110;
    rom[3394] = 25'b1111111111010110110010010;
    rom[3395] = 25'b1111111111011000010110111;
    rom[3396] = 25'b1111111111011001111011100;
    rom[3397] = 25'b1111111111011011100000000;
    rom[3398] = 25'b1111111111011101000100100;
    rom[3399] = 25'b1111111111011110101000111;
    rom[3400] = 25'b1111111111100000001101010;
    rom[3401] = 25'b1111111111100001110001011;
    rom[3402] = 25'b1111111111100011010101100;
    rom[3403] = 25'b1111111111100100111001001;
    rom[3404] = 25'b1111111111100110011100101;
    rom[3405] = 25'b1111111111100111111111111;
    rom[3406] = 25'b1111111111101001100010110;
    rom[3407] = 25'b1111111111101011000101010;
    rom[3408] = 25'b1111111111101100100111011;
    rom[3409] = 25'b1111111111101110001001001;
    rom[3410] = 25'b1111111111101111101010011;
    rom[3411] = 25'b1111111111110001001011001;
    rom[3412] = 25'b1111111111110010101011011;
    rom[3413] = 25'b1111111111110100001011001;
    rom[3414] = 25'b1111111111110101101010010;
    rom[3415] = 25'b1111111111110111001000110;
    rom[3416] = 25'b1111111111111000100110110;
    rom[3417] = 25'b1111111111111010000100000;
    rom[3418] = 25'b1111111111111011100000101;
    rom[3419] = 25'b1111111111111100111100100;
    rom[3420] = 25'b1111111111111110010111101;
    rom[3421] = 25'b1111111111111111110010000;
    rom[3422] = 25'b0000000000000001001011100;
    rom[3423] = 25'b0000000000000010100100001;
    rom[3424] = 25'b0000000000000011111100001;
    rom[3425] = 25'b0000000000000101010011001;
    rom[3426] = 25'b0000000000000110101001010;
    rom[3427] = 25'b0000000000000111111110100;
    rom[3428] = 25'b0000000000001001010010111;
    rom[3429] = 25'b0000000000001010100110001;
    rom[3430] = 25'b0000000000001011111000100;
    rom[3431] = 25'b0000000000001101001001111;
    rom[3432] = 25'b0000000000001110011010010;
    rom[3433] = 25'b0000000000001111101001100;
    rom[3434] = 25'b0000000000010000110111110;
    rom[3435] = 25'b0000000000010010000101000;
    rom[3436] = 25'b0000000000010011010001000;
    rom[3437] = 25'b0000000000010100011100000;
    rom[3438] = 25'b0000000000010101100101110;
    rom[3439] = 25'b0000000000010110101110100;
    rom[3440] = 25'b0000000000010111110110000;
    rom[3441] = 25'b0000000000011000111100010;
    rom[3442] = 25'b0000000000011010000001011;
    rom[3443] = 25'b0000000000011011000101011;
    rom[3444] = 25'b0000000000011100001000000;
    rom[3445] = 25'b0000000000011101001001101;
    rom[3446] = 25'b0000000000011110001001110;
    rom[3447] = 25'b0000000000011111001000110;
    rom[3448] = 25'b0000000000100000000110011;
    rom[3449] = 25'b0000000000100001000010111;
    rom[3450] = 25'b0000000000100001111101111;
    rom[3451] = 25'b0000000000100010110111110;
    rom[3452] = 25'b0000000000100011110000010;
    rom[3453] = 25'b0000000000100100100111011;
    rom[3454] = 25'b0000000000100101011101010;
    rom[3455] = 25'b0000000000100110010001110;
    rom[3456] = 25'b0000000000100111000100111;
    rom[3457] = 25'b0000000000100111110110110;
    rom[3458] = 25'b0000000000101000100111010;
    rom[3459] = 25'b0000000000101001010110011;
    rom[3460] = 25'b0000000000101010000100001;
    rom[3461] = 25'b0000000000101010110000100;
    rom[3462] = 25'b0000000000101011011011100;
    rom[3463] = 25'b0000000000101100000101001;
    rom[3464] = 25'b0000000000101100101101011;
    rom[3465] = 25'b0000000000101101010100001;
    rom[3466] = 25'b0000000000101101111001110;
    rom[3467] = 25'b0000000000101110011101111;
    rom[3468] = 25'b0000000000101111000000100;
    rom[3469] = 25'b0000000000101111100001111;
    rom[3470] = 25'b0000000000110000000001110;
    rom[3471] = 25'b0000000000110000100000011;
    rom[3472] = 25'b0000000000110000111101100;
    rom[3473] = 25'b0000000000110001011001010;
    rom[3474] = 25'b0000000000110001110011110;
    rom[3475] = 25'b0000000000110010001100110;
    rom[3476] = 25'b0000000000110010100100011;
    rom[3477] = 25'b0000000000110010111010110;
    rom[3478] = 25'b0000000000110011001111101;
    rom[3479] = 25'b0000000000110011100011010;
    rom[3480] = 25'b0000000000110011110101100;
    rom[3481] = 25'b0000000000110100000110011;
    rom[3482] = 25'b0000000000110100010110000;
    rom[3483] = 25'b0000000000110100100100001;
    rom[3484] = 25'b0000000000110100110001000;
    rom[3485] = 25'b0000000000110100111100100;
    rom[3486] = 25'b0000000000110101000110110;
    rom[3487] = 25'b0000000000110101001111110;
    rom[3488] = 25'b0000000000110101010111011;
    rom[3489] = 25'b0000000000110101011101110;
    rom[3490] = 25'b0000000000110101100010110;
    rom[3491] = 25'b0000000000110101100110101;
    rom[3492] = 25'b0000000000110101101001001;
    rom[3493] = 25'b0000000000110101101010011;
    rom[3494] = 25'b0000000000110101101010100;
    rom[3495] = 25'b0000000000110101101001011;
    rom[3496] = 25'b0000000000110101100111000;
    rom[3497] = 25'b0000000000110101100011011;
    rom[3498] = 25'b0000000000110101011110100;
    rom[3499] = 25'b0000000000110101011000110;
    rom[3500] = 25'b0000000000110101010001100;
    rom[3501] = 25'b0000000000110101001001010;
    rom[3502] = 25'b0000000000110100111111111;
    rom[3503] = 25'b0000000000110100110101011;
    rom[3504] = 25'b0000000000110100101001110;
    rom[3505] = 25'b0000000000110100011101000;
    rom[3506] = 25'b0000000000110100001111010;
    rom[3507] = 25'b0000000000110100000000011;
    rom[3508] = 25'b0000000000110011110000011;
    rom[3509] = 25'b0000000000110011011111011;
    rom[3510] = 25'b0000000000110011001101011;
    rom[3511] = 25'b0000000000110010111010100;
    rom[3512] = 25'b0000000000110010100110100;
    rom[3513] = 25'b0000000000110010010001101;
    rom[3514] = 25'b0000000000110001111011101;
    rom[3515] = 25'b0000000000110001100100111;
    rom[3516] = 25'b0000000000110001001101001;
    rom[3517] = 25'b0000000000110000110100011;
    rom[3518] = 25'b0000000000110000011010111;
    rom[3519] = 25'b0000000000110000000000100;
    rom[3520] = 25'b0000000000101111100101001;
    rom[3521] = 25'b0000000000101111001001000;
    rom[3522] = 25'b0000000000101110101100001;
    rom[3523] = 25'b0000000000101110001110011;
    rom[3524] = 25'b0000000000101101101111111;
    rom[3525] = 25'b0000000000101101010000100;
    rom[3526] = 25'b0000000000101100110000101;
    rom[3527] = 25'b0000000000101100001111111;
    rom[3528] = 25'b0000000000101011101110011;
    rom[3529] = 25'b0000000000101011001100010;
    rom[3530] = 25'b0000000000101010101001011;
    rom[3531] = 25'b0000000000101010000110000;
    rom[3532] = 25'b0000000000101001100001111;
    rom[3533] = 25'b0000000000101000111101001;
    rom[3534] = 25'b0000000000101000010111111;
    rom[3535] = 25'b0000000000100111110010000;
    rom[3536] = 25'b0000000000100111001011100;
    rom[3537] = 25'b0000000000100110100100101;
    rom[3538] = 25'b0000000000100101111101001;
    rom[3539] = 25'b0000000000100101010101001;
    rom[3540] = 25'b0000000000100100101100110;
    rom[3541] = 25'b0000000000100100000011110;
    rom[3542] = 25'b0000000000100011011010011;
    rom[3543] = 25'b0000000000100010110000100;
    rom[3544] = 25'b0000000000100010000110011;
    rom[3545] = 25'b0000000000100001011011110;
    rom[3546] = 25'b0000000000100000110000111;
    rom[3547] = 25'b0000000000100000000101101;
    rom[3548] = 25'b0000000000011111011010000;
    rom[3549] = 25'b0000000000011110101110000;
    rom[3550] = 25'b0000000000011110000001110;
    rom[3551] = 25'b0000000000011101010101011;
    rom[3552] = 25'b0000000000011100101000101;
    rom[3553] = 25'b0000000000011011111011100;
    rom[3554] = 25'b0000000000011011001110011;
    rom[3555] = 25'b0000000000011010100001000;
    rom[3556] = 25'b0000000000011001110011100;
    rom[3557] = 25'b0000000000011001000101101;
    rom[3558] = 25'b0000000000011000010111111;
    rom[3559] = 25'b0000000000010111101001111;
    rom[3560] = 25'b0000000000010110111011110;
    rom[3561] = 25'b0000000000010110001101100;
    rom[3562] = 25'b0000000000010101011111010;
    rom[3563] = 25'b0000000000010100110000111;
    rom[3564] = 25'b0000000000010100000010101;
    rom[3565] = 25'b0000000000010011010100001;
    rom[3566] = 25'b0000000000010010100101111;
    rom[3567] = 25'b0000000000010001110111011;
    rom[3568] = 25'b0000000000010001001001001;
    rom[3569] = 25'b0000000000010000011010111;
    rom[3570] = 25'b0000000000001111101100101;
    rom[3571] = 25'b0000000000001110111110100;
    rom[3572] = 25'b0000000000001110010000011;
    rom[3573] = 25'b0000000000001101100010100;
    rom[3574] = 25'b0000000000001100110100110;
    rom[3575] = 25'b0000000000001100000111000;
    rom[3576] = 25'b0000000000001011011001100;
    rom[3577] = 25'b0000000000001010101100001;
    rom[3578] = 25'b0000000000001001111111000;
    rom[3579] = 25'b0000000000001001010010001;
    rom[3580] = 25'b0000000000001000100101011;
    rom[3581] = 25'b0000000000000111111000110;
    rom[3582] = 25'b0000000000000111001100101;
    rom[3583] = 25'b0000000000000110100000101;
    rom[3584] = 25'b0000000000000101110100110;
    rom[3585] = 25'b0000000000000101001001011;
    rom[3586] = 25'b0000000000000100011110010;
    rom[3587] = 25'b0000000000000011110011011;
    rom[3588] = 25'b0000000000000011001000111;
    rom[3589] = 25'b0000000000000010011110110;
    rom[3590] = 25'b0000000000000001110100111;
    rom[3591] = 25'b0000000000000001001011100;
    rom[3592] = 25'b0000000000000000100010011;
    rom[3593] = 25'b1111111111111111111001110;
    rom[3594] = 25'b1111111111111111010001011;
    rom[3595] = 25'b1111111111111110101001100;
    rom[3596] = 25'b1111111111111110000010001;
    rom[3597] = 25'b1111111111111101011011000;
    rom[3598] = 25'b1111111111111100110100011;
    rom[3599] = 25'b1111111111111100001110010;
    rom[3600] = 25'b1111111111111011101000100;
    rom[3601] = 25'b1111111111111011000011010;
    rom[3602] = 25'b1111111111111010011110100;
    rom[3603] = 25'b1111111111111001111010001;
    rom[3604] = 25'b1111111111111001010110010;
    rom[3605] = 25'b1111111111111000110011000;
    rom[3606] = 25'b1111111111111000010000010;
    rom[3607] = 25'b1111111111110111101101111;
    rom[3608] = 25'b1111111111110111001100001;
    rom[3609] = 25'b1111111111110110101010111;
    rom[3610] = 25'b1111111111110110001010001;
    rom[3611] = 25'b1111111111110101101010000;
    rom[3612] = 25'b1111111111110101001010011;
    rom[3613] = 25'b1111111111110100101011011;
    rom[3614] = 25'b1111111111110100001100111;
    rom[3615] = 25'b1111111111110011101111000;
    rom[3616] = 25'b1111111111110011010001101;
    rom[3617] = 25'b1111111111110010110100111;
    rom[3618] = 25'b1111111111110010011000101;
    rom[3619] = 25'b1111111111110001111101000;
    rom[3620] = 25'b1111111111110001100010001;
    rom[3621] = 25'b1111111111110001000111110;
    rom[3622] = 25'b1111111111110000101101111;
    rom[3623] = 25'b1111111111110000010100101;
    rom[3624] = 25'b1111111111101111111100001;
    rom[3625] = 25'b1111111111101111100100001;
    rom[3626] = 25'b1111111111101111001100110;
    rom[3627] = 25'b1111111111101110110110000;
    rom[3628] = 25'b1111111111101110011111111;
    rom[3629] = 25'b1111111111101110001010011;
    rom[3630] = 25'b1111111111101101110101011;
    rom[3631] = 25'b1111111111101101100001010;
    rom[3632] = 25'b1111111111101101001101100;
    rom[3633] = 25'b1111111111101100111010100;
    rom[3634] = 25'b1111111111101100101000001;
    rom[3635] = 25'b1111111111101100010110011;
    rom[3636] = 25'b1111111111101100000101010;
    rom[3637] = 25'b1111111111101011110100110;
    rom[3638] = 25'b1111111111101011100100111;
    rom[3639] = 25'b1111111111101011010101101;
    rom[3640] = 25'b1111111111101011000111000;
    rom[3641] = 25'b1111111111101010111001000;
    rom[3642] = 25'b1111111111101010101011101;
    rom[3643] = 25'b1111111111101010011110111;
    rom[3644] = 25'b1111111111101010010010110;
    rom[3645] = 25'b1111111111101010000111010;
    rom[3646] = 25'b1111111111101001111100011;
    rom[3647] = 25'b1111111111101001110010001;
    rom[3648] = 25'b1111111111101001101000011;
    rom[3649] = 25'b1111111111101001011111011;
    rom[3650] = 25'b1111111111101001010110111;
    rom[3651] = 25'b1111111111101001001111000;
    rom[3652] = 25'b1111111111101001000111111;
    rom[3653] = 25'b1111111111101001000001010;
    rom[3654] = 25'b1111111111101000111011010;
    rom[3655] = 25'b1111111111101000110101110;
    rom[3656] = 25'b1111111111101000110001000;
    rom[3657] = 25'b1111111111101000101100101;
    rom[3658] = 25'b1111111111101000101000111;
    rom[3659] = 25'b1111111111101000100101111;
    rom[3660] = 25'b1111111111101000100011011;
    rom[3661] = 25'b1111111111101000100001010;
    rom[3662] = 25'b1111111111101000011111111;
    rom[3663] = 25'b1111111111101000011111000;
    rom[3664] = 25'b1111111111101000011110110;
    rom[3665] = 25'b1111111111101000011111000;
    rom[3666] = 25'b1111111111101000011111110;
    rom[3667] = 25'b1111111111101000100001001;
    rom[3668] = 25'b1111111111101000100011000;
    rom[3669] = 25'b1111111111101000100101010;
    rom[3670] = 25'b1111111111101000101000010;
    rom[3671] = 25'b1111111111101000101011100;
    rom[3672] = 25'b1111111111101000101111100;
    rom[3673] = 25'b1111111111101000110011111;
    rom[3674] = 25'b1111111111101000111000110;
    rom[3675] = 25'b1111111111101000111110001;
    rom[3676] = 25'b1111111111101001000100000;
    rom[3677] = 25'b1111111111101001001010010;
    rom[3678] = 25'b1111111111101001010001001;
    rom[3679] = 25'b1111111111101001011000010;
    rom[3680] = 25'b1111111111101001100000000;
    rom[3681] = 25'b1111111111101001101000001;
    rom[3682] = 25'b1111111111101001110000110;
    rom[3683] = 25'b1111111111101001111001101;
    rom[3684] = 25'b1111111111101010000011001;
    rom[3685] = 25'b1111111111101010001101000;
    rom[3686] = 25'b1111111111101010010111001;
    rom[3687] = 25'b1111111111101010100001110;
    rom[3688] = 25'b1111111111101010101100111;
    rom[3689] = 25'b1111111111101010111000010;
    rom[3690] = 25'b1111111111101011000100000;
    rom[3691] = 25'b1111111111101011010000001;
    rom[3692] = 25'b1111111111101011011100100;
    rom[3693] = 25'b1111111111101011101001011;
    rom[3694] = 25'b1111111111101011110110101;
    rom[3695] = 25'b1111111111101100000100001;
    rom[3696] = 25'b1111111111101100010001111;
    rom[3697] = 25'b1111111111101100100000000;
    rom[3698] = 25'b1111111111101100101110100;
    rom[3699] = 25'b1111111111101100111101010;
    rom[3700] = 25'b1111111111101101001100010;
    rom[3701] = 25'b1111111111101101011011101;
    rom[3702] = 25'b1111111111101101101011001;
    rom[3703] = 25'b1111111111101101111011000;
    rom[3704] = 25'b1111111111101110001011001;
    rom[3705] = 25'b1111111111101110011011100;
    rom[3706] = 25'b1111111111101110101100000;
    rom[3707] = 25'b1111111111101110111100111;
    rom[3708] = 25'b1111111111101111001110000;
    rom[3709] = 25'b1111111111101111011111010;
    rom[3710] = 25'b1111111111101111110000101;
    rom[3711] = 25'b1111111111110000000010010;
    rom[3712] = 25'b1111111111110000010100001;
    rom[3713] = 25'b1111111111110000100110001;
    rom[3714] = 25'b1111111111110000111000011;
    rom[3715] = 25'b1111111111110001001010110;
    rom[3716] = 25'b1111111111110001011101010;
    rom[3717] = 25'b1111111111110001101111111;
    rom[3718] = 25'b1111111111110010000010101;
    rom[3719] = 25'b1111111111110010010101101;
    rom[3720] = 25'b1111111111110010101000101;
    rom[3721] = 25'b1111111111110010111011110;
    rom[3722] = 25'b1111111111110011001111000;
    rom[3723] = 25'b1111111111110011100010011;
    rom[3724] = 25'b1111111111110011110101110;
    rom[3725] = 25'b1111111111110100001001010;
    rom[3726] = 25'b1111111111110100011100111;
    rom[3727] = 25'b1111111111110100110000100;
    rom[3728] = 25'b1111111111110101000100010;
    rom[3729] = 25'b1111111111110101010111111;
    rom[3730] = 25'b1111111111110101101011110;
    rom[3731] = 25'b1111111111110101111111100;
    rom[3732] = 25'b1111111111110110010011011;
    rom[3733] = 25'b1111111111110110100111010;
    rom[3734] = 25'b1111111111110110111011001;
    rom[3735] = 25'b1111111111110111001111000;
    rom[3736] = 25'b1111111111110111100010111;
    rom[3737] = 25'b1111111111110111110110101;
    rom[3738] = 25'b1111111111111000001010100;
    rom[3739] = 25'b1111111111111000011110010;
    rom[3740] = 25'b1111111111111000110010000;
    rom[3741] = 25'b1111111111111001000101110;
    rom[3742] = 25'b1111111111111001011001100;
    rom[3743] = 25'b1111111111111001101101000;
    rom[3744] = 25'b1111111111111010000000101;
    rom[3745] = 25'b1111111111111010010100001;
    rom[3746] = 25'b1111111111111010100111101;
    rom[3747] = 25'b1111111111111010111010111;
    rom[3748] = 25'b1111111111111011001110001;
    rom[3749] = 25'b1111111111111011100001010;
    rom[3750] = 25'b1111111111111011110100011;
    rom[3751] = 25'b1111111111111100000111010;
    rom[3752] = 25'b1111111111111100011010001;
    rom[3753] = 25'b1111111111111100101100110;
    rom[3754] = 25'b1111111111111100111111011;
    rom[3755] = 25'b1111111111111101010001110;
    rom[3756] = 25'b1111111111111101100100001;
    rom[3757] = 25'b1111111111111101110110011;
    rom[3758] = 25'b1111111111111110001000011;
    rom[3759] = 25'b1111111111111110011010010;
    rom[3760] = 25'b1111111111111110101100000;
    rom[3761] = 25'b1111111111111110111101101;
    rom[3762] = 25'b1111111111111111001111000;
    rom[3763] = 25'b1111111111111111100000010;
    rom[3764] = 25'b1111111111111111110001010;
    rom[3765] = 25'b0000000000000000000010001;
    rom[3766] = 25'b0000000000000000010010110;
    rom[3767] = 25'b0000000000000000100011010;
    rom[3768] = 25'b0000000000000000110011101;
    rom[3769] = 25'b0000000000000001000011110;
    rom[3770] = 25'b0000000000000001010011101;
    rom[3771] = 25'b0000000000000001100011011;
    rom[3772] = 25'b0000000000000001110010111;
    rom[3773] = 25'b0000000000000010000010001;
    rom[3774] = 25'b0000000000000010010001010;
    rom[3775] = 25'b0000000000000010100000001;
    rom[3776] = 25'b0000000000000010101110110;
    rom[3777] = 25'b0000000000000010111101001;
    rom[3778] = 25'b0000000000000011001011011;
    rom[3779] = 25'b0000000000000011011001011;
    rom[3780] = 25'b0000000000000011100111000;
    rom[3781] = 25'b0000000000000011110100100;
    rom[3782] = 25'b0000000000000100000001110;
    rom[3783] = 25'b0000000000000100001110111;
    rom[3784] = 25'b0000000000000100011011101;
    rom[3785] = 25'b0000000000000100101000001;
    rom[3786] = 25'b0000000000000100110100011;
    rom[3787] = 25'b0000000000000101000000011;
    rom[3788] = 25'b0000000000000101001100010;
    rom[3789] = 25'b0000000000000101010111110;
    rom[3790] = 25'b0000000000000101100011000;
    rom[3791] = 25'b0000000000000101101110001;
    rom[3792] = 25'b0000000000000101111000110;
    rom[3793] = 25'b0000000000000110000011011;
    rom[3794] = 25'b0000000000000110001101101;
    rom[3795] = 25'b0000000000000110010111101;
    rom[3796] = 25'b0000000000000110100001010;
    rom[3797] = 25'b0000000000000110101010110;
    rom[3798] = 25'b0000000000000110110100000;
    rom[3799] = 25'b0000000000000110111101000;
    rom[3800] = 25'b0000000000000111000101101;
    rom[3801] = 25'b0000000000000111001110000;
    rom[3802] = 25'b0000000000000111010110001;
    rom[3803] = 25'b0000000000000111011110000;
    rom[3804] = 25'b0000000000000111100101110;
    rom[3805] = 25'b0000000000000111101101000;
    rom[3806] = 25'b0000000000000111110100001;
    rom[3807] = 25'b0000000000000111111011000;
    rom[3808] = 25'b0000000000001000000001100;
    rom[3809] = 25'b0000000000001000000111110;
    rom[3810] = 25'b0000000000001000001101111;
    rom[3811] = 25'b0000000000001000010011101;
    rom[3812] = 25'b0000000000001000011001001;
    rom[3813] = 25'b0000000000001000011110100;
    rom[3814] = 25'b0000000000001000100011011;
    rom[3815] = 25'b0000000000001000101000001;
    rom[3816] = 25'b0000000000001000101100101;
    rom[3817] = 25'b0000000000001000110000111;
    rom[3818] = 25'b0000000000001000110100111;
    rom[3819] = 25'b0000000000001000111000100;
    rom[3820] = 25'b0000000000001000111100001;
    rom[3821] = 25'b0000000000001000111111010;
    rom[3822] = 25'b0000000000001001000010010;
    rom[3823] = 25'b0000000000001001000101000;
    rom[3824] = 25'b0000000000001001000111100;
    rom[3825] = 25'b0000000000001001001001110;
    rom[3826] = 25'b0000000000001001001011101;
    rom[3827] = 25'b0000000000001001001101100;
    rom[3828] = 25'b0000000000001001001111000;
    rom[3829] = 25'b0000000000001001010000010;
    rom[3830] = 25'b0000000000001001010001011;
    rom[3831] = 25'b0000000000001001010010010;
    rom[3832] = 25'b0000000000001001010010110;
    rom[3833] = 25'b0000000000001001010011001;
    rom[3834] = 25'b0000000000001001010011010;
    rom[3835] = 25'b0000000000001001010011010;
    rom[3836] = 25'b0000000000001001010010111;
    rom[3837] = 25'b0000000000001001010010011;
    rom[3838] = 25'b0000000000001001010001101;
    rom[3839] = 25'b0000000000001001010000110;
    rom[3840] = 25'b0000000000001001001111101;
    rom[3841] = 25'b0000000000001001001110010;
    rom[3842] = 25'b0000000000001001001100110;
    rom[3843] = 25'b0000000000001001001010111;
    rom[3844] = 25'b0000000000001001001001000;
    rom[3845] = 25'b0000000000001001000110111;
    rom[3846] = 25'b0000000000001001000100101;
    rom[3847] = 25'b0000000000001001000010001;
    rom[3848] = 25'b0000000000001000111111011;
    rom[3849] = 25'b0000000000001000111100100;
    rom[3850] = 25'b0000000000001000111001011;
    rom[3851] = 25'b0000000000001000110110010;
    rom[3852] = 25'b0000000000001000110010111;
    rom[3853] = 25'b0000000000001000101111010;
    rom[3854] = 25'b0000000000001000101011100;
    rom[3855] = 25'b0000000000001000100111101;
    rom[3856] = 25'b0000000000001000100011101;
    rom[3857] = 25'b0000000000001000011111100;
    rom[3858] = 25'b0000000000001000011011001;
    rom[3859] = 25'b0000000000001000010110101;
    rom[3860] = 25'b0000000000001000010010000;
    rom[3861] = 25'b0000000000001000001101010;
    rom[3862] = 25'b0000000000001000001000010;
    rom[3863] = 25'b0000000000001000000011010;
    rom[3864] = 25'b0000000000000111111110001;
    rom[3865] = 25'b0000000000000111111000110;
    rom[3866] = 25'b0000000000000111110011011;
    rom[3867] = 25'b0000000000000111101101111;
    rom[3868] = 25'b0000000000000111101000010;
    rom[3869] = 25'b0000000000000111100010100;
    rom[3870] = 25'b0000000000000111011100101;
    rom[3871] = 25'b0000000000000111010110101;
    rom[3872] = 25'b0000000000000111010000101;
    rom[3873] = 25'b0000000000000111001010100;
    rom[3874] = 25'b0000000000000111000100010;
    rom[3875] = 25'b0000000000000110111101111;
    rom[3876] = 25'b0000000000000110110111100;
    rom[3877] = 25'b0000000000000110110000111;
    rom[3878] = 25'b0000000000000110101010011;
    rom[3879] = 25'b0000000000000110100011110;
    rom[3880] = 25'b0000000000000110011101000;
    rom[3881] = 25'b0000000000000110010110001;
    rom[3882] = 25'b0000000000000110001111011;
    rom[3883] = 25'b0000000000000110001000100;
    rom[3884] = 25'b0000000000000110000001100;
    rom[3885] = 25'b0000000000000101111010011;
    rom[3886] = 25'b0000000000000101110011010;
    rom[3887] = 25'b0000000000000101101100010;
    rom[3888] = 25'b0000000000000101100101000;
    rom[3889] = 25'b0000000000000101011101111;
    rom[3890] = 25'b0000000000000101010110101;
    rom[3891] = 25'b0000000000000101001111011;
    rom[3892] = 25'b0000000000000101001000000;
    rom[3893] = 25'b0000000000000101000000110;
    rom[3894] = 25'b0000000000000100111001011;
    rom[3895] = 25'b0000000000000100110010000;
    rom[3896] = 25'b0000000000000100101010110;
    rom[3897] = 25'b0000000000000100100011010;
    rom[3898] = 25'b0000000000000100011011111;
    rom[3899] = 25'b0000000000000100010100011;
    rom[3900] = 25'b0000000000000100001101000;
    rom[3901] = 25'b0000000000000100000101101;
    rom[3902] = 25'b0000000000000011111110010;
    rom[3903] = 25'b0000000000000011110110110;
    rom[3904] = 25'b0000000000000011101111011;
    rom[3905] = 25'b0000000000000011101000000;
    rom[3906] = 25'b0000000000000011100000101;
    rom[3907] = 25'b0000000000000011011001011;
    rom[3908] = 25'b0000000000000011010010000;
    rom[3909] = 25'b0000000000000011001010101;
    rom[3910] = 25'b0000000000000011000011011;
    rom[3911] = 25'b0000000000000010111100001;
    rom[3912] = 25'b0000000000000010110101000;
    rom[3913] = 25'b0000000000000010101101110;
    rom[3914] = 25'b0000000000000010100110101;
    rom[3915] = 25'b0000000000000010011111100;
    rom[3916] = 25'b0000000000000010011000100;
    rom[3917] = 25'b0000000000000010010001011;
    rom[3918] = 25'b0000000000000010001010100;
    rom[3919] = 25'b0000000000000010000011100;
    rom[3920] = 25'b0000000000000001111100101;
    rom[3921] = 25'b0000000000000001110101110;
    rom[3922] = 25'b0000000000000001101111000;
    rom[3923] = 25'b0000000000000001101000010;
    rom[3924] = 25'b0000000000000001100001101;
    rom[3925] = 25'b0000000000000001011011000;
    rom[3926] = 25'b0000000000000001010100100;
    rom[3927] = 25'b0000000000000001001110000;
    rom[3928] = 25'b0000000000000001000111101;
    rom[3929] = 25'b0000000000000001000001010;
    rom[3930] = 25'b0000000000000000111011000;
    rom[3931] = 25'b0000000000000000110100111;
    rom[3932] = 25'b0000000000000000101110110;
    rom[3933] = 25'b0000000000000000101000101;
    rom[3934] = 25'b0000000000000000100010110;
    rom[3935] = 25'b0000000000000000011100111;
    rom[3936] = 25'b0000000000000000010111000;
    rom[3937] = 25'b0000000000000000010001011;
    rom[3938] = 25'b0000000000000000001011101;
    rom[3939] = 25'b0000000000000000000110001;
    rom[3940] = 25'b0000000000000000000000101;
    rom[3941] = 25'b1111111111111111111011011;
    rom[3942] = 25'b1111111111111111110110000;
    rom[3943] = 25'b1111111111111111110000111;
    rom[3944] = 25'b1111111111111111101011110;
    rom[3945] = 25'b1111111111111111100110101;
    rom[3946] = 25'b1111111111111111100001110;
    rom[3947] = 25'b1111111111111111011100111;
    rom[3948] = 25'b1111111111111111011000001;
    rom[3949] = 25'b1111111111111111010011100;
    rom[3950] = 25'b1111111111111111001110111;
    rom[3951] = 25'b1111111111111111001010011;
    rom[3952] = 25'b1111111111111111000110001;
    rom[3953] = 25'b1111111111111111000001111;
    rom[3954] = 25'b1111111111111110111101101;
    rom[3955] = 25'b1111111111111110111001100;
    rom[3956] = 25'b1111111111111110110101100;
    rom[3957] = 25'b1111111111111110110001101;
    rom[3958] = 25'b1111111111111110101101111;
    rom[3959] = 25'b1111111111111110101010001;
    rom[3960] = 25'b1111111111111110100110100;
    rom[3961] = 25'b1111111111111110100011001;
    rom[3962] = 25'b1111111111111110011111101;
    rom[3963] = 25'b1111111111111110011100011;
    rom[3964] = 25'b1111111111111110011001010;
    rom[3965] = 25'b1111111111111110010110000;
    rom[3966] = 25'b1111111111111110010011000;
    rom[3967] = 25'b1111111111111110010000001;
    rom[3968] = 25'b1111111111111110001101011;
    rom[3969] = 25'b1111111111111110001010101;
    rom[3970] = 25'b1111111111111110001000000;
    rom[3971] = 25'b1111111111111110000101100;
    rom[3972] = 25'b1111111111111110000011000;
    rom[3973] = 25'b1111111111111110000000110;
    rom[3974] = 25'b1111111111111101111110100;
    rom[3975] = 25'b1111111111111101111100011;
    rom[3976] = 25'b1111111111111101111010011;
    rom[3977] = 25'b1111111111111101111000011;
    rom[3978] = 25'b1111111111111101110110100;
    rom[3979] = 25'b1111111111111101110100110;
    rom[3980] = 25'b1111111111111101110011001;
    rom[3981] = 25'b1111111111111101110001100;
    rom[3982] = 25'b1111111111111101110000000;
    rom[3983] = 25'b1111111111111101101110101;
    rom[3984] = 25'b1111111111111101101101010;
    rom[3985] = 25'b1111111111111101101100001;
    rom[3986] = 25'b1111111111111101101011000;
    rom[3987] = 25'b1111111111111101101001111;
    rom[3988] = 25'b1111111111111101101000111;
    rom[3989] = 25'b1111111111111101101000001;
    rom[3990] = 25'b1111111111111101100111010;
    rom[3991] = 25'b1111111111111101100110100;
    rom[3992] = 25'b1111111111111101100101111;
    rom[3993] = 25'b1111111111111101100101010;
    rom[3994] = 25'b1111111111111101100100111;
    rom[3995] = 25'b1111111111111101100100100;
    rom[3996] = 25'b1111111111111101100100001;
    rom[3997] = 25'b1111111111111101100011111;
    rom[3998] = 25'b1111111111111101100011110;
    rom[3999] = 25'b1111111111111101100011100;
    rom[4000] = 25'b1111111111111101100011100;
    rom[4001] = 25'b1111111111111101100011100;
    rom[4002] = 25'b1111111111111101100011101;
    rom[4003] = 25'b1111111111111101100011110;
    rom[4004] = 25'b1111111111111101100100001;
    rom[4005] = 25'b1111111111111101100100011;
    rom[4006] = 25'b1111111111111101100100101;
    rom[4007] = 25'b1111111111111101100101001;
    rom[4008] = 25'b1111111111111101100101101;
    rom[4009] = 25'b1111111111111101100110000;
    rom[4010] = 25'b1111111111111101100110110;
    rom[4011] = 25'b1111111111111101100111011;
    rom[4012] = 25'b1111111111111101101000000;
    rom[4013] = 25'b1111111111111101101000110;
    rom[4014] = 25'b1111111111111101101001100;
    rom[4015] = 25'b1111111111111101101010011;
    rom[4016] = 25'b1111111111111101101011010;
    rom[4017] = 25'b1111111111111101101100010;
    rom[4018] = 25'b1111111111111101101101001;
    rom[4019] = 25'b1111111111111101101110001;
    rom[4020] = 25'b1111111111111101101111001;
    rom[4021] = 25'b1111111111111101110000010;
    rom[4022] = 25'b1111111111111101110001011;
    rom[4023] = 25'b1111111111111101110010100;
    rom[4024] = 25'b1111111111111101110011110;
    rom[4025] = 25'b1111111111111101110101000;
    rom[4026] = 25'b1111111111111101110110010;
    rom[4027] = 25'b1111111111111101110111100;
    rom[4028] = 25'b1111111111111101111000111;
    rom[4029] = 25'b1111111111111101111010001;
    rom[4030] = 25'b1111111111111101111011101;
    rom[4031] = 25'b1111111111111101111100111;
    rom[4032] = 25'b1111111111111101111110010;
    rom[4033] = 25'b1111111111111101111111101;
    rom[4034] = 25'b1111111111111110000001001;
    rom[4035] = 25'b1111111111111110000010100;
    rom[4036] = 25'b1111111111111110000100000;
    rom[4037] = 25'b1111111111111110000101100;
    rom[4038] = 25'b1111111111111110000111000;
    rom[4039] = 25'b1111111111111110001000100;
    rom[4040] = 25'b1111111111111110001010000;
    rom[4041] = 25'b1111111111111110001011100;
    rom[4042] = 25'b1111111111111110001101000;
    rom[4043] = 25'b1111111111111110001110100;
    rom[4044] = 25'b1111111111111110010000001;
    rom[4045] = 25'b1111111111111110010001101;
    rom[4046] = 25'b1111111111111110010011000;
    rom[4047] = 25'b1111111111111110010100100;
    rom[4048] = 25'b1111111111111110010110000;
    rom[4049] = 25'b1111111111111110010111100;
    rom[4050] = 25'b1111111111111110011001000;
    rom[4051] = 25'b1111111111111110011010100;
    rom[4052] = 25'b1111111111111110011100000;
    rom[4053] = 25'b1111111111111110011101011;
    rom[4054] = 25'b1111111111111110011110111;
    rom[4055] = 25'b1111111111111110100000010;
    rom[4056] = 25'b1111111111111110100001110;
    rom[4057] = 25'b1111111111111110100011001;
    rom[4058] = 25'b1111111111111110100100100;
    rom[4059] = 25'b1111111111111110100101110;
    rom[4060] = 25'b1111111111111110100111010;
    rom[4061] = 25'b1111111111111110101000100;
    rom[4062] = 25'b1111111111111110101001110;
    rom[4063] = 25'b1111111111111110101011000;
    rom[4064] = 25'b1111111111111110101100011;
    rom[4065] = 25'b1111111111111110101101100;
    rom[4066] = 25'b1111111111111110101110101;
    rom[4067] = 25'b1111111111111110101111111;
    rom[4068] = 25'b1111111111111110110001000;
    rom[4069] = 25'b1111111111111110110010000;
    rom[4070] = 25'b1111111111111110110011001;
    rom[4071] = 25'b1111111111111110110100001;
    rom[4072] = 25'b1111111111111110110101001;
    rom[4073] = 25'b1111111111111110110110001;
    rom[4074] = 25'b1111111111111110110111000;
    rom[4075] = 25'b1111111111111110110111111;
    rom[4076] = 25'b1111111111111110111000111;
    rom[4077] = 25'b1111111111111110111001100;
    rom[4078] = 25'b1111111111111110111010011;
    rom[4079] = 25'b1111111111111110111011001;
    rom[4080] = 25'b1111111111111110111011110;
    rom[4081] = 25'b1111111111111110111100100;
    rom[4082] = 25'b1111111111111110111101001;
    rom[4083] = 25'b1111111111111110111101101;
    rom[4084] = 25'b1111111111111110111110010;
    rom[4085] = 25'b1111111111111110111110110;
    rom[4086] = 25'b1111111111111110111111001;
    rom[4087] = 25'b1111111111111110111111101;
    rom[4088] = 25'b1111111111111111000000000;
    rom[4089] = 25'b1111111111111111000000010;
    rom[4090] = 25'b1111111111111111000000100;
    rom[4091] = 25'b1111111111111111000000111;
    rom[4092] = 25'b1111111111111111000001000;
    rom[4093] = 25'b1111111111111111000001010;
    rom[4094] = 25'b1111111111111111000001010;
    rom[4095] = 25'b1111111111111111000001011;
end

// port a
always @(posedge clk)
begin
    if (wea_d == 1'b1) begin
      rom[addra_d] <= dia_d;
    end
    wea_d <= wea;
    dia_d <= dia;
    addra_d <= addra;
end

// port b
always @(posedge clk)
begin
    addrb_d <= addrb;
    rom_pipea <= rom[addrb_d];
    dob_d <= rom_pipea;
end

endmodule
