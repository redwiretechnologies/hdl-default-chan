// SPDX-License-Identifier: Apache-2.0

// Tags are 7-bits wide.

localparam CHAN_TAG_FIRST = 'd07;
