// Tags are 7-bits wide.

localparam CHAN_TAG_FIRST = 'd07;
