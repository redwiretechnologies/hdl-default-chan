//
// Macros used only in Simulation
//
//
`ifndef SIM_BIN_WRITE
//`define SIM_BIN_WRITE 1
`endif
