// SPDX-License-Identifier: Apache-2.0

/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : cic_M256_N1_R1_iw5_0_correction_sp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data
//
//
/*****************************************************************************/


module cic_M256_N1_R1_iw5_0_correction_sp_rom
(
  input clk,

  input [8:0] addra,
  output [12:0] doa
);

(* rom_style = "block" *) reg [12:0] rom [511:0];
reg [8:0] addra_d;
reg [12:0] doa_d;
reg [12:0] rom_pipea;

assign doa = doa_d;

initial
begin
    rom[0] = 13'b0000100000000;
    rom[1] = 13'b0000100000000;
    rom[2] = 13'b0000010000000;
    rom[3] = 13'b0000001010101;
    rom[4] = 13'b0000001000000;
    rom[5] = 13'b0000000110011;
    rom[6] = 13'b0000000101011;
    rom[7] = 13'b0000000100101;
    rom[8] = 13'b0000000100000;
    rom[9] = 13'b0000000011100;
    rom[10] = 13'b0000000011010;
    rom[11] = 13'b0000000010111;
    rom[12] = 13'b0000000010101;
    rom[13] = 13'b0000000010100;
    rom[14] = 13'b0000000010010;
    rom[15] = 13'b0000000010001;
    rom[16] = 13'b0000000010000;
    rom[17] = 13'b0000000001111;
    rom[18] = 13'b0000000001110;
    rom[19] = 13'b0000000001101;
    rom[20] = 13'b0000000001101;
    rom[21] = 13'b0000000001100;
    rom[22] = 13'b0000000001100;
    rom[23] = 13'b0000000001011;
    rom[24] = 13'b0000000001011;
    rom[25] = 13'b0000000001010;
    rom[26] = 13'b0000000001010;
    rom[27] = 13'b0000000001001;
    rom[28] = 13'b0000000001001;
    rom[29] = 13'b0000000001001;
    rom[30] = 13'b0000000001001;
    rom[31] = 13'b0000000001000;
    rom[32] = 13'b0000000001000;
    rom[33] = 13'b0000000001000;
    rom[34] = 13'b0000000001000;
    rom[35] = 13'b0000000000111;
    rom[36] = 13'b0000000000111;
    rom[37] = 13'b0000000000111;
    rom[38] = 13'b0000000000111;
    rom[39] = 13'b0000000000111;
    rom[40] = 13'b0000000000110;
    rom[41] = 13'b0000000000110;
    rom[42] = 13'b0000000000110;
    rom[43] = 13'b0000000000110;
    rom[44] = 13'b0000000000110;
    rom[45] = 13'b0000000000110;
    rom[46] = 13'b0000000000110;
    rom[47] = 13'b0000000000101;
    rom[48] = 13'b0000000000101;
    rom[49] = 13'b0000000000101;
    rom[50] = 13'b0000000000101;
    rom[51] = 13'b0000000000101;
    rom[52] = 13'b0000000000101;
    rom[53] = 13'b0000000000101;
    rom[54] = 13'b0000000000101;
    rom[55] = 13'b0000000000101;
    rom[56] = 13'b0000000000101;
    rom[57] = 13'b0000000000100;
    rom[58] = 13'b0000000000100;
    rom[59] = 13'b0000000000100;
    rom[60] = 13'b0000000000100;
    rom[61] = 13'b0000000000100;
    rom[62] = 13'b0000000000100;
    rom[63] = 13'b0000000000100;
    rom[64] = 13'b0000000000100;
    rom[65] = 13'b0000000000100;
    rom[66] = 13'b0000000000100;
    rom[67] = 13'b0000000000100;
    rom[68] = 13'b0000000000100;
    rom[69] = 13'b0000000000100;
    rom[70] = 13'b0000000000100;
    rom[71] = 13'b0000000000100;
    rom[72] = 13'b0000000000100;
    rom[73] = 13'b0000000000100;
    rom[74] = 13'b0000000000011;
    rom[75] = 13'b0000000000011;
    rom[76] = 13'b0000000000011;
    rom[77] = 13'b0000000000011;
    rom[78] = 13'b0000000000011;
    rom[79] = 13'b0000000000011;
    rom[80] = 13'b0000000000011;
    rom[81] = 13'b0000000000011;
    rom[82] = 13'b0000000000011;
    rom[83] = 13'b0000000000011;
    rom[84] = 13'b0000000000011;
    rom[85] = 13'b0000000000011;
    rom[86] = 13'b0000000000011;
    rom[87] = 13'b0000000000011;
    rom[88] = 13'b0000000000011;
    rom[89] = 13'b0000000000011;
    rom[90] = 13'b0000000000011;
    rom[91] = 13'b0000000000011;
    rom[92] = 13'b0000000000011;
    rom[93] = 13'b0000000000011;
    rom[94] = 13'b0000000000011;
    rom[95] = 13'b0000000000011;
    rom[96] = 13'b0000000000011;
    rom[97] = 13'b0000000000011;
    rom[98] = 13'b0000000000011;
    rom[99] = 13'b0000000000011;
    rom[100] = 13'b0000000000011;
    rom[101] = 13'b0000000000011;
    rom[102] = 13'b0000000000011;
    rom[103] = 13'b0000000000010;
    rom[104] = 13'b0000000000010;
    rom[105] = 13'b0000000000010;
    rom[106] = 13'b0000000000010;
    rom[107] = 13'b0000000000010;
    rom[108] = 13'b0000000000010;
    rom[109] = 13'b0000000000010;
    rom[110] = 13'b0000000000010;
    rom[111] = 13'b0000000000010;
    rom[112] = 13'b0000000000010;
    rom[113] = 13'b0000000000010;
    rom[114] = 13'b0000000000010;
    rom[115] = 13'b0000000000010;
    rom[116] = 13'b0000000000010;
    rom[117] = 13'b0000000000010;
    rom[118] = 13'b0000000000010;
    rom[119] = 13'b0000000000010;
    rom[120] = 13'b0000000000010;
    rom[121] = 13'b0000000000010;
    rom[122] = 13'b0000000000010;
    rom[123] = 13'b0000000000010;
    rom[124] = 13'b0000000000010;
    rom[125] = 13'b0000000000010;
    rom[126] = 13'b0000000000010;
    rom[127] = 13'b0000000000010;
    rom[128] = 13'b0000000000010;
    rom[129] = 13'b0000000000010;
    rom[130] = 13'b0000000000010;
    rom[131] = 13'b0000000000010;
    rom[132] = 13'b0000000000010;
    rom[133] = 13'b0000000000010;
    rom[134] = 13'b0000000000010;
    rom[135] = 13'b0000000000010;
    rom[136] = 13'b0000000000010;
    rom[137] = 13'b0000000000010;
    rom[138] = 13'b0000000000010;
    rom[139] = 13'b0000000000010;
    rom[140] = 13'b0000000000010;
    rom[141] = 13'b0000000000010;
    rom[142] = 13'b0000000000010;
    rom[143] = 13'b0000000000010;
    rom[144] = 13'b0000000000010;
    rom[145] = 13'b0000000000010;
    rom[146] = 13'b0000000000010;
    rom[147] = 13'b0000000000010;
    rom[148] = 13'b0000000000010;
    rom[149] = 13'b0000000000010;
    rom[150] = 13'b0000000000010;
    rom[151] = 13'b0000000000010;
    rom[152] = 13'b0000000000010;
    rom[153] = 13'b0000000000010;
    rom[154] = 13'b0000000000010;
    rom[155] = 13'b0000000000010;
    rom[156] = 13'b0000000000010;
    rom[157] = 13'b0000000000010;
    rom[158] = 13'b0000000000010;
    rom[159] = 13'b0000000000010;
    rom[160] = 13'b0000000000010;
    rom[161] = 13'b0000000000010;
    rom[162] = 13'b0000000000010;
    rom[163] = 13'b0000000000010;
    rom[164] = 13'b0000000000010;
    rom[165] = 13'b0000000000010;
    rom[166] = 13'b0000000000010;
    rom[167] = 13'b0000000000010;
    rom[168] = 13'b0000000000010;
    rom[169] = 13'b0000000000010;
    rom[170] = 13'b0000000000010;
    rom[171] = 13'b0000000000001;
    rom[172] = 13'b0000000000001;
    rom[173] = 13'b0000000000001;
    rom[174] = 13'b0000000000001;
    rom[175] = 13'b0000000000001;
    rom[176] = 13'b0000000000001;
    rom[177] = 13'b0000000000001;
    rom[178] = 13'b0000000000001;
    rom[179] = 13'b0000000000001;
    rom[180] = 13'b0000000000001;
    rom[181] = 13'b0000000000001;
    rom[182] = 13'b0000000000001;
    rom[183] = 13'b0000000000001;
    rom[184] = 13'b0000000000001;
    rom[185] = 13'b0000000000001;
    rom[186] = 13'b0000000000001;
    rom[187] = 13'b0000000000001;
    rom[188] = 13'b0000000000001;
    rom[189] = 13'b0000000000001;
    rom[190] = 13'b0000000000001;
    rom[191] = 13'b0000000000001;
    rom[192] = 13'b0000000000001;
    rom[193] = 13'b0000000000001;
    rom[194] = 13'b0000000000001;
    rom[195] = 13'b0000000000001;
    rom[196] = 13'b0000000000001;
    rom[197] = 13'b0000000000001;
    rom[198] = 13'b0000000000001;
    rom[199] = 13'b0000000000001;
    rom[200] = 13'b0000000000001;
    rom[201] = 13'b0000000000001;
    rom[202] = 13'b0000000000001;
    rom[203] = 13'b0000000000001;
    rom[204] = 13'b0000000000001;
    rom[205] = 13'b0000000000001;
    rom[206] = 13'b0000000000001;
    rom[207] = 13'b0000000000001;
    rom[208] = 13'b0000000000001;
    rom[209] = 13'b0000000000001;
    rom[210] = 13'b0000000000001;
    rom[211] = 13'b0000000000001;
    rom[212] = 13'b0000000000001;
    rom[213] = 13'b0000000000001;
    rom[214] = 13'b0000000000001;
    rom[215] = 13'b0000000000001;
    rom[216] = 13'b0000000000001;
    rom[217] = 13'b0000000000001;
    rom[218] = 13'b0000000000001;
    rom[219] = 13'b0000000000001;
    rom[220] = 13'b0000000000001;
    rom[221] = 13'b0000000000001;
    rom[222] = 13'b0000000000001;
    rom[223] = 13'b0000000000001;
    rom[224] = 13'b0000000000001;
    rom[225] = 13'b0000000000001;
    rom[226] = 13'b0000000000001;
    rom[227] = 13'b0000000000001;
    rom[228] = 13'b0000000000001;
    rom[229] = 13'b0000000000001;
    rom[230] = 13'b0000000000001;
    rom[231] = 13'b0000000000001;
    rom[232] = 13'b0000000000001;
    rom[233] = 13'b0000000000001;
    rom[234] = 13'b0000000000001;
    rom[235] = 13'b0000000000001;
    rom[236] = 13'b0000000000001;
    rom[237] = 13'b0000000000001;
    rom[238] = 13'b0000000000001;
    rom[239] = 13'b0000000000001;
    rom[240] = 13'b0000000000001;
    rom[241] = 13'b0000000000001;
    rom[242] = 13'b0000000000001;
    rom[243] = 13'b0000000000001;
    rom[244] = 13'b0000000000001;
    rom[245] = 13'b0000000000001;
    rom[246] = 13'b0000000000001;
    rom[247] = 13'b0000000000001;
    rom[248] = 13'b0000000000001;
    rom[249] = 13'b0000000000001;
    rom[250] = 13'b0000000000001;
    rom[251] = 13'b0000000000001;
    rom[252] = 13'b0000000000001;
    rom[253] = 13'b0000000000001;
    rom[254] = 13'b0000000000001;
    rom[255] = 13'b0000000000001;
    rom[256] = 13'b0000000000001;
    rom[257] = 13'b0000000000000;
    rom[258] = 13'b0000000000000;
    rom[259] = 13'b0000000000000;
    rom[260] = 13'b0000000000000;
    rom[261] = 13'b0000000000000;
    rom[262] = 13'b0000000000000;
    rom[263] = 13'b0000000000000;
    rom[264] = 13'b0000000000000;
    rom[265] = 13'b0000000000000;
    rom[266] = 13'b0000000000000;
    rom[267] = 13'b0000000000000;
    rom[268] = 13'b0000000000000;
    rom[269] = 13'b0000000000000;
    rom[270] = 13'b0000000000000;
    rom[271] = 13'b0000000000000;
    rom[272] = 13'b0000000000000;
    rom[273] = 13'b0000000000000;
    rom[274] = 13'b0000000000000;
    rom[275] = 13'b0000000000000;
    rom[276] = 13'b0000000000000;
    rom[277] = 13'b0000000000000;
    rom[278] = 13'b0000000000000;
    rom[279] = 13'b0000000000000;
    rom[280] = 13'b0000000000000;
    rom[281] = 13'b0000000000000;
    rom[282] = 13'b0000000000000;
    rom[283] = 13'b0000000000000;
    rom[284] = 13'b0000000000000;
    rom[285] = 13'b0000000000000;
    rom[286] = 13'b0000000000000;
    rom[287] = 13'b0000000000000;
    rom[288] = 13'b0000000000000;
    rom[289] = 13'b0000000000000;
    rom[290] = 13'b0000000000000;
    rom[291] = 13'b0000000000000;
    rom[292] = 13'b0000000000000;
    rom[293] = 13'b0000000000000;
    rom[294] = 13'b0000000000000;
    rom[295] = 13'b0000000000000;
    rom[296] = 13'b0000000000000;
    rom[297] = 13'b0000000000000;
    rom[298] = 13'b0000000000000;
    rom[299] = 13'b0000000000000;
    rom[300] = 13'b0000000000000;
    rom[301] = 13'b0000000000000;
    rom[302] = 13'b0000000000000;
    rom[303] = 13'b0000000000000;
    rom[304] = 13'b0000000000000;
    rom[305] = 13'b0000000000000;
    rom[306] = 13'b0000000000000;
    rom[307] = 13'b0000000000000;
    rom[308] = 13'b0000000000000;
    rom[309] = 13'b0000000000000;
    rom[310] = 13'b0000000000000;
    rom[311] = 13'b0000000000000;
    rom[312] = 13'b0000000000000;
    rom[313] = 13'b0000000000000;
    rom[314] = 13'b0000000000000;
    rom[315] = 13'b0000000000000;
    rom[316] = 13'b0000000000000;
    rom[317] = 13'b0000000000000;
    rom[318] = 13'b0000000000000;
    rom[319] = 13'b0000000000000;
    rom[320] = 13'b0000000000000;
    rom[321] = 13'b0000000000000;
    rom[322] = 13'b0000000000000;
    rom[323] = 13'b0000000000000;
    rom[324] = 13'b0000000000000;
    rom[325] = 13'b0000000000000;
    rom[326] = 13'b0000000000000;
    rom[327] = 13'b0000000000000;
    rom[328] = 13'b0000000000000;
    rom[329] = 13'b0000000000000;
    rom[330] = 13'b0000000000000;
    rom[331] = 13'b0000000000000;
    rom[332] = 13'b0000000000000;
    rom[333] = 13'b0000000000000;
    rom[334] = 13'b0000000000000;
    rom[335] = 13'b0000000000000;
    rom[336] = 13'b0000000000000;
    rom[337] = 13'b0000000000000;
    rom[338] = 13'b0000000000000;
    rom[339] = 13'b0000000000000;
    rom[340] = 13'b0000000000000;
    rom[341] = 13'b0000000000000;
    rom[342] = 13'b0000000000000;
    rom[343] = 13'b0000000000000;
    rom[344] = 13'b0000000000000;
    rom[345] = 13'b0000000000000;
    rom[346] = 13'b0000000000000;
    rom[347] = 13'b0000000000000;
    rom[348] = 13'b0000000000000;
    rom[349] = 13'b0000000000000;
    rom[350] = 13'b0000000000000;
    rom[351] = 13'b0000000000000;
    rom[352] = 13'b0000000000000;
    rom[353] = 13'b0000000000000;
    rom[354] = 13'b0000000000000;
    rom[355] = 13'b0000000000000;
    rom[356] = 13'b0000000000000;
    rom[357] = 13'b0000000000000;
    rom[358] = 13'b0000000000000;
    rom[359] = 13'b0000000000000;
    rom[360] = 13'b0000000000000;
    rom[361] = 13'b0000000000000;
    rom[362] = 13'b0000000000000;
    rom[363] = 13'b0000000000000;
    rom[364] = 13'b0000000000000;
    rom[365] = 13'b0000000000000;
    rom[366] = 13'b0000000000000;
    rom[367] = 13'b0000000000000;
    rom[368] = 13'b0000000000000;
    rom[369] = 13'b0000000000000;
    rom[370] = 13'b0000000000000;
    rom[371] = 13'b0000000000000;
    rom[372] = 13'b0000000000000;
    rom[373] = 13'b0000000000000;
    rom[374] = 13'b0000000000000;
    rom[375] = 13'b0000000000000;
    rom[376] = 13'b0000000000000;
    rom[377] = 13'b0000000000000;
    rom[378] = 13'b0000000000000;
    rom[379] = 13'b0000000000000;
    rom[380] = 13'b0000000000000;
    rom[381] = 13'b0000000000000;
    rom[382] = 13'b0000000000000;
    rom[383] = 13'b0000000000000;
    rom[384] = 13'b0000000000000;
    rom[385] = 13'b0000000000000;
    rom[386] = 13'b0000000000000;
    rom[387] = 13'b0000000000000;
    rom[388] = 13'b0000000000000;
    rom[389] = 13'b0000000000000;
    rom[390] = 13'b0000000000000;
    rom[391] = 13'b0000000000000;
    rom[392] = 13'b0000000000000;
    rom[393] = 13'b0000000000000;
    rom[394] = 13'b0000000000000;
    rom[395] = 13'b0000000000000;
    rom[396] = 13'b0000000000000;
    rom[397] = 13'b0000000000000;
    rom[398] = 13'b0000000000000;
    rom[399] = 13'b0000000000000;
    rom[400] = 13'b0000000000000;
    rom[401] = 13'b0000000000000;
    rom[402] = 13'b0000000000000;
    rom[403] = 13'b0000000000000;
    rom[404] = 13'b0000000000000;
    rom[405] = 13'b0000000000000;
    rom[406] = 13'b0000000000000;
    rom[407] = 13'b0000000000000;
    rom[408] = 13'b0000000000000;
    rom[409] = 13'b0000000000000;
    rom[410] = 13'b0000000000000;
    rom[411] = 13'b0000000000000;
    rom[412] = 13'b0000000000000;
    rom[413] = 13'b0000000000000;
    rom[414] = 13'b0000000000000;
    rom[415] = 13'b0000000000000;
    rom[416] = 13'b0000000000000;
    rom[417] = 13'b0000000000000;
    rom[418] = 13'b0000000000000;
    rom[419] = 13'b0000000000000;
    rom[420] = 13'b0000000000000;
    rom[421] = 13'b0000000000000;
    rom[422] = 13'b0000000000000;
    rom[423] = 13'b0000000000000;
    rom[424] = 13'b0000000000000;
    rom[425] = 13'b0000000000000;
    rom[426] = 13'b0000000000000;
    rom[427] = 13'b0000000000000;
    rom[428] = 13'b0000000000000;
    rom[429] = 13'b0000000000000;
    rom[430] = 13'b0000000000000;
    rom[431] = 13'b0000000000000;
    rom[432] = 13'b0000000000000;
    rom[433] = 13'b0000000000000;
    rom[434] = 13'b0000000000000;
    rom[435] = 13'b0000000000000;
    rom[436] = 13'b0000000000000;
    rom[437] = 13'b0000000000000;
    rom[438] = 13'b0000000000000;
    rom[439] = 13'b0000000000000;
    rom[440] = 13'b0000000000000;
    rom[441] = 13'b0000000000000;
    rom[442] = 13'b0000000000000;
    rom[443] = 13'b0000000000000;
    rom[444] = 13'b0000000000000;
    rom[445] = 13'b0000000000000;
    rom[446] = 13'b0000000000000;
    rom[447] = 13'b0000000000000;
    rom[448] = 13'b0000000000000;
    rom[449] = 13'b0000000000000;
    rom[450] = 13'b0000000000000;
    rom[451] = 13'b0000000000000;
    rom[452] = 13'b0000000000000;
    rom[453] = 13'b0000000000000;
    rom[454] = 13'b0000000000000;
    rom[455] = 13'b0000000000000;
    rom[456] = 13'b0000000000000;
    rom[457] = 13'b0000000000000;
    rom[458] = 13'b0000000000000;
    rom[459] = 13'b0000000000000;
    rom[460] = 13'b0000000000000;
    rom[461] = 13'b0000000000000;
    rom[462] = 13'b0000000000000;
    rom[463] = 13'b0000000000000;
    rom[464] = 13'b0000000000000;
    rom[465] = 13'b0000000000000;
    rom[466] = 13'b0000000000000;
    rom[467] = 13'b0000000000000;
    rom[468] = 13'b0000000000000;
    rom[469] = 13'b0000000000000;
    rom[470] = 13'b0000000000000;
    rom[471] = 13'b0000000000000;
    rom[472] = 13'b0000000000000;
    rom[473] = 13'b0000000000000;
    rom[474] = 13'b0000000000000;
    rom[475] = 13'b0000000000000;
    rom[476] = 13'b0000000000000;
    rom[477] = 13'b0000000000000;
    rom[478] = 13'b0000000000000;
    rom[479] = 13'b0000000000000;
    rom[480] = 13'b0000000000000;
    rom[481] = 13'b0000000000000;
    rom[482] = 13'b0000000000000;
    rom[483] = 13'b0000000000000;
    rom[484] = 13'b0000000000000;
    rom[485] = 13'b0000000000000;
    rom[486] = 13'b0000000000000;
    rom[487] = 13'b0000000000000;
    rom[488] = 13'b0000000000000;
    rom[489] = 13'b0000000000000;
    rom[490] = 13'b0000000000000;
    rom[491] = 13'b0000000000000;
    rom[492] = 13'b0000000000000;
    rom[493] = 13'b0000000000000;
    rom[494] = 13'b0000000000000;
    rom[495] = 13'b0000000000000;
    rom[496] = 13'b0000000000000;
    rom[497] = 13'b0000000000000;
    rom[498] = 13'b0000000000000;
    rom[499] = 13'b0000000000000;
    rom[500] = 13'b0000000000000;
    rom[501] = 13'b0000000000000;
    rom[502] = 13'b0000000000000;
    rom[503] = 13'b0000000000000;
    rom[504] = 13'b0000000000000;
    rom[505] = 13'b0000000000000;
    rom[506] = 13'b0000000000000;
    rom[507] = 13'b0000000000000;
    rom[508] = 13'b0000000000000;
    rom[509] = 13'b0000000000000;
    rom[510] = 13'b0000000000000;
    rom[511] = 13'b0000000000000;
end

// port a
always @(posedge clk)
begin
    addra_d <= addra;
    rom_pipea <= rom[addra_d];
    doa_d <= rom_pipea;
end

endmodule
